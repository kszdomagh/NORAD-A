//////////////////////////////////////////////////////////////////////////////
/*
 Module name:   ending_screen_rom
 Author:        kszdom
 Description:   ROM memory for ending screen


  _   _ _    _  _____ _      ______          _____                        
 | \ | | |  | |/ ____| |    |  ____|   /\   |  __ \                       
 |  \| | |  | | |    | |    | |__     /  \  | |__) |                      
 | . ` | |  | | |    | |    |  __|   / /\ \ |  _  /                       
 | |\  | |__| | |____| |____| |____ / ____ \| | \ \                       
 |_| \_|\____/_\_____|______|______/_/_ __\_\_|__\_\  _____   ____  _   _ 
     /\   |  __ \|  \/  |   /\   / ____|  ____|  __ \|  __ \ / __ \| \ | |
    /  \  | |__) | \  / |  /  \ | |  __| |__  | |  | | |  | | |  | |  \| |
   / /\ \ |  _  /| |\/| | / /\ \| | |_ |  __| | |  | | |  | | |  | | . ` |
  / ____ \| | \ \| |  | |/ ____ \ |__| | |____| |__| | |__| | |__| | |\  |
 /_/___ \_\_|_ \_\_| _|_/_/__  \_\_____|______|_____/|_____/ \____/|_| \_|
 |_   _|/ ____| | \ | |  ____|   /\   |  __ \                             
   | | | (___   |  \| | |__     /  \  | |__) |                            
   | |  \___ \  | . ` |  __|   / /\ \ |  _  /                             
  _| |_ ____) | | |\  | |____ / ____ \| | \ \                             
 |_____|_____/  |_| \_|______/_/    \_\_|  \_\ 

 */
//////////////////////////////////////////////////////////////////////////////



module end_screen_rom #(
    parameter int ADDRESSWIDTH = 4,  // 4 bits => 16 entries
    parameter int DATAWIDTH = 18  // 8+8+1+1 = 18 bits
)(
    input logic [ADDRESSWIDTH-1:0] addr,
    output logic [DATAWIDTH-1:0] data_out
);

    always_comb begin
        unique case (addr)
            //                  x       y       line    pos

            0: data_out = {8'd54, 8'd187, 1'b0, 1'b1};
            1: data_out = {8'd69, 8'd187, 1'b1, 1'b0};
            2: data_out = {8'd69, 8'd194, 1'b1, 1'b0};
            3: data_out = {8'd54, 8'd194, 1'b1, 1'b0};
            4: data_out = {8'd54, 8'd187, 1'b1, 1'b0};
            5: data_out = {8'd46, 8'd163, 1'b0, 1'b1};
            6: data_out = {8'd53, 8'd163, 1'b1, 1'b0};
            7: data_out = {8'd53, 8'd186, 1'b1, 1'b0};
            8: data_out = {8'd46, 8'd186, 1'b1, 1'b0};
            9: data_out = {8'd46, 8'd163, 1'b1, 1'b0};
            10: data_out = {8'd54, 8'd155, 1'b0, 1'b1};
            11: data_out = {8'd69, 8'd155, 1'b1, 1'b0};
            12: data_out = {8'd69, 8'd162, 1'b1, 1'b0};
            13: data_out = {8'd54, 8'd162, 1'b1, 1'b0};
            14: data_out = {8'd54, 8'd155, 1'b1, 1'b0};
            15: data_out = {8'd62, 8'd171, 1'b0, 1'b1};
            16: data_out = {8'd77, 8'd171, 1'b1, 1'b0};
            17: data_out = {8'd77, 8'd178, 1'b1, 1'b0};
            18: data_out = {8'd62, 8'd178, 1'b1, 1'b0};
            19: data_out = {8'd62, 8'd171, 1'b1, 1'b0};
            20: data_out = {8'd70, 8'd171, 1'b0, 1'b1};
            21: data_out = {8'd70, 8'd163, 1'b1, 1'b0};
            22: data_out = {8'd77, 8'd163, 1'b1, 1'b0};
            23: data_out = {8'd77, 8'd171, 1'b1, 1'b0};
            24: data_out = {8'd86, 8'd155, 1'b0, 1'b1};
            25: data_out = {8'd93, 8'd155, 1'b1, 1'b0};
            26: data_out = {8'd93, 8'd186, 1'b1, 1'b0};
            27: data_out = {8'd86, 8'd186, 1'b1, 1'b0};
            28: data_out = {8'd86, 8'd155, 1'b1, 1'b0};
            29: data_out = {8'd94, 8'd187, 1'b0, 1'b1};
            30: data_out = {8'd109, 8'd187, 1'b1, 1'b0};
            31: data_out = {8'd109, 8'd194, 1'b1, 1'b0};
            32: data_out = {8'd94, 8'd194, 1'b1, 1'b0};
            33: data_out = {8'd94, 8'd187, 1'b1, 1'b0};
            34: data_out = {8'd110, 8'd155, 1'b0, 1'b1};
            35: data_out = {8'd117, 8'd155, 1'b1, 1'b0};
            36: data_out = {8'd117, 8'd186, 1'b1, 1'b0};
            37: data_out = {8'd110, 8'd186, 1'b1, 1'b0};
            38: data_out = {8'd110, 8'd155, 1'b1, 1'b0};
            39: data_out = {8'd93, 8'd171, 1'b0, 1'b1};
            40: data_out = {8'd110, 8'd171, 1'b1, 1'b0};
            41: data_out = {8'd93, 8'd178, 1'b0, 1'b1};
            42: data_out = {8'd110, 8'd178, 1'b1, 1'b0};
            43: data_out = {8'd126, 8'd155, 1'b0, 1'b1};
            44: data_out = {8'd133, 8'd155, 1'b1, 1'b0};
            45: data_out = {8'd133, 8'd194, 1'b1, 1'b0};
            46: data_out = {8'd126, 8'd194, 1'b1, 1'b0};
            47: data_out = {8'd126, 8'd155, 1'b1, 1'b0};
            48: data_out = {8'd142, 8'd171, 1'b0, 1'b1};
            49: data_out = {8'd149, 8'd171, 1'b1, 1'b0};
            50: data_out = {8'd149, 8'd178, 1'b1, 1'b0};
            51: data_out = {8'd142, 8'd178, 1'b1, 1'b0};
            52: data_out = {8'd142, 8'd171, 1'b1, 1'b0};
            53: data_out = {8'd158, 8'd155, 1'b0, 1'b1};
            54: data_out = {8'd165, 8'd155, 1'b1, 1'b0};
            55: data_out = {8'd165, 8'd194, 1'b1, 1'b0};
            56: data_out = {8'd158, 8'd194, 1'b1, 1'b0};
            57: data_out = {8'd158, 8'd155, 1'b1, 1'b0};
            58: data_out = {8'd133, 8'd179, 1'b0, 1'b1};
            59: data_out = {8'd141, 8'd179, 1'b1, 1'b0};
            60: data_out = {8'd141, 8'd186, 1'b1, 1'b0};
            61: data_out = {8'd133, 8'd186, 1'b1, 1'b0};
            62: data_out = {8'd158, 8'd179, 1'b0, 1'b1};
            63: data_out = {8'd150, 8'd179, 1'b1, 1'b0};
            64: data_out = {8'd150, 8'd186, 1'b1, 1'b0};
            65: data_out = {8'd158, 8'd186, 1'b1, 1'b0};
            66: data_out = {8'd174, 8'd155, 1'b0, 1'b1};
            67: data_out = {8'd181, 8'd155, 1'b1, 1'b0};
            68: data_out = {8'd181, 8'd194, 1'b1, 1'b0};
            69: data_out = {8'd174, 8'd194, 1'b1, 1'b0};
            70: data_out = {8'd174, 8'd155, 1'b1, 1'b0};
            71: data_out = {8'd181, 8'd155, 1'b0, 1'b1};
            72: data_out = {8'd205, 8'd155, 1'b1, 1'b0};
            73: data_out = {8'd205, 8'd162, 1'b1, 1'b0};
            74: data_out = {8'd181, 8'd162, 1'b1, 1'b0};
            75: data_out = {8'd181, 8'd171, 1'b0, 1'b1};
            76: data_out = {8'd197, 8'd171, 1'b1, 1'b0};
            77: data_out = {8'd197, 8'd178, 1'b1, 1'b0};
            78: data_out = {8'd181, 8'd178, 1'b1, 1'b0};
            79: data_out = {8'd181, 8'd187, 1'b0, 1'b1};
            80: data_out = {8'd205, 8'd187, 1'b1, 1'b0};
            81: data_out = {8'd205, 8'd194, 1'b1, 1'b0};
            82: data_out = {8'd181, 8'd194, 1'b1, 1'b0};
            83: data_out = {8'd47, 8'd83, 1'b0, 1'b1};
            84: data_out = {8'd54, 8'd83, 1'b1, 1'b0};
            85: data_out = {8'd54, 8'd106, 1'b1, 1'b0};
            86: data_out = {8'd47, 8'd106, 1'b1, 1'b0};
            87: data_out = {8'd47, 8'd83, 1'b1, 1'b0};
            88: data_out = {8'd55, 8'd75, 1'b0, 1'b1};
            89: data_out = {8'd70, 8'd75, 1'b1, 1'b0};
            90: data_out = {8'd70, 8'd82, 1'b1, 1'b0};
            91: data_out = {8'd55, 8'd82, 1'b1, 1'b0};
            92: data_out = {8'd55, 8'd75, 1'b1, 1'b0};
            93: data_out = {8'd71, 8'd83, 1'b0, 1'b1};
            94: data_out = {8'd78, 8'd83, 1'b1, 1'b0};
            95: data_out = {8'd78, 8'd106, 1'b1, 1'b0};
            96: data_out = {8'd71, 8'd106, 1'b1, 1'b0};
            97: data_out = {8'd71, 8'd83, 1'b1, 1'b0};
            98: data_out = {8'd55, 8'd107, 1'b0, 1'b1};
            99: data_out = {8'd70, 8'd107, 1'b1, 1'b0};
            100: data_out = {8'd70, 8'd114, 1'b1, 1'b0};
            101: data_out = {8'd55, 8'd114, 1'b1, 1'b0};
            102: data_out = {8'd55, 8'd107, 1'b1, 1'b0};
            103: data_out = {8'd87, 8'd99, 1'b0, 1'b1};
            104: data_out = {8'd94, 8'd99, 1'b1, 1'b0};
            105: data_out = {8'd94, 8'd114, 1'b1, 1'b0};
            106: data_out = {8'd87, 8'd114, 1'b1, 1'b0};
            107: data_out = {8'd87, 8'd99, 1'b1, 1'b0};
            108: data_out = {8'd95, 8'd83, 1'b0, 1'b1};
            109: data_out = {8'd102, 8'd83, 1'b1, 1'b0};
            110: data_out = {8'd102, 8'd98, 1'b1, 1'b0};
            111: data_out = {8'd95, 8'd98, 1'b1, 1'b0};
            112: data_out = {8'd95, 8'd83, 1'b1, 1'b0};
            113: data_out = {8'd103, 8'd75, 1'b0, 1'b1};
            114: data_out = {8'd110, 8'd75, 1'b1, 1'b0};
            115: data_out = {8'd110, 8'd82, 1'b1, 1'b0};
            116: data_out = {8'd103, 8'd82, 1'b1, 1'b0};
            117: data_out = {8'd103, 8'd75, 1'b1, 1'b0};
            118: data_out = {8'd111, 8'd83, 1'b0, 1'b1};
            119: data_out = {8'd118, 8'd83, 1'b1, 1'b0};
            120: data_out = {8'd118, 8'd98, 1'b1, 1'b0};
            121: data_out = {8'd111, 8'd98, 1'b1, 1'b0};
            122: data_out = {8'd111, 8'd83, 1'b1, 1'b0};
            123: data_out = {8'd119, 8'd99, 1'b0, 1'b1};
            124: data_out = {8'd126, 8'd99, 1'b1, 1'b0};
            125: data_out = {8'd126, 8'd114, 1'b1, 1'b0};
            126: data_out = {8'd119, 8'd114, 1'b1, 1'b0};
            127: data_out = {8'd119, 8'd99, 1'b1, 1'b0};
            128: data_out = {8'd135, 8'd75, 1'b0, 1'b1};
            129: data_out = {8'd142, 8'd75, 1'b1, 1'b0};
            130: data_out = {8'd142, 8'd114, 1'b1, 1'b0};
            131: data_out = {8'd135, 8'd114, 1'b1, 1'b0};
            132: data_out = {8'd135, 8'd75, 1'b1, 1'b0};
            133: data_out = {8'd142, 8'd75, 1'b0, 1'b1};
            134: data_out = {8'd166, 8'd75, 1'b1, 1'b0};
            135: data_out = {8'd166, 8'd82, 1'b1, 1'b0};
            136: data_out = {8'd142, 8'd82, 1'b1, 1'b0};
            137: data_out = {8'd142, 8'd91, 1'b0, 1'b1};
            138: data_out = {8'd158, 8'd91, 1'b1, 1'b0};
            139: data_out = {8'd158, 8'd98, 1'b1, 1'b0};
            140: data_out = {8'd142, 8'd98, 1'b1, 1'b0};
            141: data_out = {8'd142, 8'd107, 1'b0, 1'b1};
            142: data_out = {8'd166, 8'd107, 1'b1, 1'b0};
            143: data_out = {8'd166, 8'd114, 1'b1, 1'b0};
            144: data_out = {8'd142, 8'd114, 1'b1, 1'b0};
            145: data_out = {8'd175, 8'd74, 1'b0, 1'b1};
            146: data_out = {8'd182, 8'd74, 1'b1, 1'b0};
            147: data_out = {8'd182, 8'd114, 1'b1, 1'b0};
            148: data_out = {8'd175, 8'd114, 1'b1, 1'b0};
            149: data_out = {8'd175, 8'd74, 1'b1, 1'b0};
            150: data_out = {8'd199, 8'd99, 1'b0, 1'b1};
            151: data_out = {8'd206, 8'd99, 1'b1, 1'b0};
            152: data_out = {8'd206, 8'd106, 1'b1, 1'b0};
            153: data_out = {8'd199, 8'd106, 1'b1, 1'b0};
            154: data_out = {8'd199, 8'd99, 1'b1, 1'b0};
            155: data_out = {8'd199, 8'd75, 1'b0, 1'b1};
            156: data_out = {8'd206, 8'd75, 1'b1, 1'b0};
            157: data_out = {8'd206, 8'd82, 1'b1, 1'b0};
            158: data_out = {8'd199, 8'd82, 1'b1, 1'b0};
            159: data_out = {8'd199, 8'd75, 1'b1, 1'b0};
            160: data_out = {8'd182, 8'd107, 1'b0, 1'b1};
            161: data_out = {8'd198, 8'd107, 1'b1, 1'b0};
            162: data_out = {8'd198, 8'd114, 1'b1, 1'b0};
            163: data_out = {8'd182, 8'd114, 1'b1, 1'b0};
            164: data_out = {8'd182, 8'd91, 1'b0, 1'b1};
            165: data_out = {8'd198, 8'd91, 1'b1, 1'b0};
            166: data_out = {8'd198, 8'd98, 1'b1, 1'b0};
            167: data_out = {8'd182, 8'd98, 1'b1, 1'b0};
            168: data_out = {8'd191, 8'd91, 1'b0, 1'b1};
            169: data_out = {8'd191, 8'd83, 1'b1, 1'b0};
            170: data_out = {8'd198, 8'd83, 1'b1, 1'b0};
            171: data_out = {8'd198, 8'd91, 1'b1, 1'b0};
            172: data_out = {8'd198, 8'd91, 1'b1, 1'b1};    // RESET



            default: data_out = '0;
        endcase
    end

endmodule
