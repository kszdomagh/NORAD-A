//////////////////////////////////////////////////////////////////////////////
/*
 Module name:   uwu_rom
 Author:        kszdom
 Description:   test ROM image module 


  _   _ _    _  _____ _      ______          _____                        
 | \ | | |  | |/ ____| |    |  ____|   /\   |  __ \                       
 |  \| | |  | | |    | |    | |__     /  \  | |__) |                      
 | . ` | |  | | |    | |    |  __|   / /\ \ |  _  /                       
 | |\  | |__| | |____| |____| |____ / ____ \| | \ \                       
 |_| \_|\____/_\_____|______|______/_/_ __\_\_|__\_\  _____   ____  _   _ 
     /\   |  __ \|  \/  |   /\   / ____|  ____|  __ \|  __ \ / __ \| \ | |
    /  \  | |__) | \  / |  /  \ | |  __| |__  | |  | | |  | | |  | |  \| |
   / /\ \ |  _  /| |\/| | / /\ \| | |_ |  __| | |  | | |  | | |  | | . ` |
  / ____ \| | \ \| |  | |/ ____ \ |__| | |____| |__| | |__| | |__| | |\  |
 /_/___ \_\_|_ \_\_| _|_/_/__  \_\_____|______|_____/|_____/ \____/|_| \_|
 |_   _|/ ____| | \ | |  ____|   /\   |  __ \                             
   | | | (___   |  \| | |__     /  \  | |__) |                            
   | |  \___ \  | . ` |  __|   / /\ \ |  _  /                             
  _| |_ ____) | | |\  | |____ / ____ \| | \ \                             
 |_____|_____/  |_| \_|______/_/    \_\_|  \_\ 

 */
//////////////////////////////////////////////////////////////////////////////



module start_rom #(
    parameter int ADDRESSWIDTH = 16,  // 4 bits => 16 entries
    parameter int DATAWIDTH = 18  // 8+8+1+1 = 18 bits
)(
    input logic [ADDRESSWIDTH-1:0] addr,
    output logic [DATAWIDTH-1:0] data_out
);


    always_comb begin
        unique case (addr)


0: data_out = {8'd146, 8'd7, 1'b1, 1'b0};
1: data_out = {8'd147, 8'd7, 1'b1, 1'b0};
2: data_out = {8'd148, 8'd7, 1'b1, 1'b0};
3: data_out = {8'd149, 8'd7, 1'b1, 1'b0};
4: data_out = {8'd150, 8'd7, 1'b1, 1'b0};
5: data_out = {8'd151, 8'd7, 1'b1, 1'b0};
6: data_out = {8'd146, 8'd8, 1'b1, 1'b0};
7: data_out = {8'd147, 8'd8, 1'b1, 1'b0};
8: data_out = {8'd148, 8'd8, 1'b1, 1'b0};
9: data_out = {8'd149, 8'd8, 1'b1, 1'b0};
10: data_out = {8'd150, 8'd8, 1'b1, 1'b0};
11: data_out = {8'd151, 8'd8, 1'b1, 1'b0};
12: data_out = {8'd146, 8'd9, 1'b1, 1'b0};
13: data_out = {8'd147, 8'd9, 1'b1, 1'b0};
14: data_out = {8'd148, 8'd9, 1'b1, 1'b0};
15: data_out = {8'd149, 8'd9, 1'b1, 1'b0};
16: data_out = {8'd150, 8'd9, 1'b1, 1'b0};
17: data_out = {8'd151, 8'd9, 1'b1, 1'b0};
18: data_out = {8'd146, 8'd10, 1'b1, 1'b0};
19: data_out = {8'd147, 8'd10, 1'b1, 1'b0};
20: data_out = {8'd148, 8'd10, 1'b1, 1'b0};
21: data_out = {8'd149, 8'd10, 1'b1, 1'b0};
22: data_out = {8'd150, 8'd10, 1'b1, 1'b0};
23: data_out = {8'd151, 8'd10, 1'b1, 1'b0};
24: data_out = {8'd146, 8'd11, 1'b1, 1'b0};
25: data_out = {8'd147, 8'd11, 1'b1, 1'b0};
26: data_out = {8'd148, 8'd11, 1'b1, 1'b0};
27: data_out = {8'd149, 8'd11, 1'b1, 1'b0};
28: data_out = {8'd150, 8'd11, 1'b1, 1'b0};
29: data_out = {8'd151, 8'd11, 1'b1, 1'b0};
30: data_out = {8'd146, 8'd12, 1'b1, 1'b0};
31: data_out = {8'd147, 8'd12, 1'b1, 1'b0};
32: data_out = {8'd148, 8'd12, 1'b1, 1'b0};
33: data_out = {8'd149, 8'd12, 1'b1, 1'b0};
34: data_out = {8'd150, 8'd12, 1'b1, 1'b0};
35: data_out = {8'd151, 8'd12, 1'b1, 1'b0};
36: data_out = {8'd146, 8'd13, 1'b1, 1'b0};
37: data_out = {8'd147, 8'd13, 1'b1, 1'b0};
38: data_out = {8'd148, 8'd13, 1'b1, 1'b0};
39: data_out = {8'd149, 8'd13, 1'b1, 1'b0};
40: data_out = {8'd150, 8'd13, 1'b1, 1'b0};
41: data_out = {8'd151, 8'd13, 1'b1, 1'b0};
42: data_out = {8'd146, 8'd14, 1'b1, 1'b0};
43: data_out = {8'd147, 8'd14, 1'b1, 1'b0};
44: data_out = {8'd148, 8'd14, 1'b1, 1'b0};
45: data_out = {8'd149, 8'd14, 1'b1, 1'b0};
46: data_out = {8'd150, 8'd14, 1'b1, 1'b0};
47: data_out = {8'd151, 8'd14, 1'b1, 1'b0};
48: data_out = {8'd146, 8'd15, 1'b1, 1'b0};
49: data_out = {8'd147, 8'd15, 1'b1, 1'b0};
50: data_out = {8'd148, 8'd15, 1'b1, 1'b0};
51: data_out = {8'd149, 8'd15, 1'b1, 1'b0};
52: data_out = {8'd150, 8'd15, 1'b1, 1'b0};
53: data_out = {8'd151, 8'd15, 1'b1, 1'b0};
54: data_out = {8'd146, 8'd16, 1'b1, 1'b0};
55: data_out = {8'd147, 8'd16, 1'b1, 1'b0};
56: data_out = {8'd148, 8'd16, 1'b1, 1'b0};
57: data_out = {8'd149, 8'd16, 1'b1, 1'b0};
58: data_out = {8'd150, 8'd16, 1'b1, 1'b0};
59: data_out = {8'd151, 8'd16, 1'b1, 1'b0};
60: data_out = {8'd146, 8'd17, 1'b1, 1'b0};
61: data_out = {8'd147, 8'd17, 1'b1, 1'b0};
62: data_out = {8'd148, 8'd17, 1'b1, 1'b0};
63: data_out = {8'd149, 8'd17, 1'b1, 1'b0};
64: data_out = {8'd150, 8'd17, 1'b1, 1'b0};
65: data_out = {8'd151, 8'd17, 1'b1, 1'b0};
66: data_out = {8'd146, 8'd18, 1'b1, 1'b0};
67: data_out = {8'd147, 8'd18, 1'b1, 1'b0};
68: data_out = {8'd148, 8'd18, 1'b1, 1'b0};
69: data_out = {8'd149, 8'd18, 1'b1, 1'b0};
70: data_out = {8'd150, 8'd18, 1'b1, 1'b0};
71: data_out = {8'd151, 8'd18, 1'b1, 1'b0};
72: data_out = {8'd146, 8'd19, 1'b1, 1'b0};
73: data_out = {8'd147, 8'd19, 1'b1, 1'b0};
74: data_out = {8'd148, 8'd19, 1'b1, 1'b0};
75: data_out = {8'd149, 8'd19, 1'b1, 1'b0};
76: data_out = {8'd150, 8'd19, 1'b1, 1'b0};
77: data_out = {8'd151, 8'd19, 1'b1, 1'b0};
78: data_out = {8'd8, 8'd20, 1'b1, 1'b0};
79: data_out = {8'd9, 8'd20, 1'b1, 1'b0};
80: data_out = {8'd10, 8'd20, 1'b1, 1'b0};
81: data_out = {8'd11, 8'd20, 1'b1, 1'b0};
82: data_out = {8'd12, 8'd20, 1'b1, 1'b0};
83: data_out = {8'd13, 8'd20, 1'b1, 1'b0};
84: data_out = {8'd14, 8'd20, 1'b1, 1'b0};
85: data_out = {8'd15, 8'd20, 1'b1, 1'b0};
86: data_out = {8'd16, 8'd20, 1'b1, 1'b0};
87: data_out = {8'd17, 8'd20, 1'b1, 1'b0};
88: data_out = {8'd18, 8'd20, 1'b1, 1'b0};
89: data_out = {8'd19, 8'd20, 1'b1, 1'b0};
90: data_out = {8'd20, 8'd20, 1'b1, 1'b0};
91: data_out = {8'd21, 8'd20, 1'b1, 1'b0};
92: data_out = {8'd22, 8'd20, 1'b1, 1'b0};
93: data_out = {8'd23, 8'd20, 1'b1, 1'b0};
94: data_out = {8'd24, 8'd20, 1'b1, 1'b0};
95: data_out = {8'd25, 8'd20, 1'b1, 1'b0};
96: data_out = {8'd26, 8'd20, 1'b1, 1'b0};
97: data_out = {8'd27, 8'd20, 1'b1, 1'b0};
98: data_out = {8'd28, 8'd20, 1'b1, 1'b0};
99: data_out = {8'd38, 8'd20, 1'b1, 1'b0};
100: data_out = {8'd39, 8'd20, 1'b1, 1'b0};
101: data_out = {8'd40, 8'd20, 1'b1, 1'b0};
102: data_out = {8'd41, 8'd20, 1'b1, 1'b0};
103: data_out = {8'd42, 8'd20, 1'b1, 1'b0};
104: data_out = {8'd43, 8'd20, 1'b1, 1'b0};
105: data_out = {8'd44, 8'd20, 1'b1, 1'b0};
106: data_out = {8'd45, 8'd20, 1'b1, 1'b0};
107: data_out = {8'd46, 8'd20, 1'b1, 1'b0};
108: data_out = {8'd47, 8'd20, 1'b1, 1'b0};
109: data_out = {8'd48, 8'd20, 1'b1, 1'b0};
110: data_out = {8'd49, 8'd20, 1'b1, 1'b0};
111: data_out = {8'd50, 8'd20, 1'b1, 1'b0};
112: data_out = {8'd51, 8'd20, 1'b1, 1'b0};
113: data_out = {8'd52, 8'd20, 1'b1, 1'b0};
114: data_out = {8'd53, 8'd20, 1'b1, 1'b0};
115: data_out = {8'd54, 8'd20, 1'b1, 1'b0};
116: data_out = {8'd55, 8'd20, 1'b1, 1'b0};
117: data_out = {8'd56, 8'd20, 1'b1, 1'b0};
118: data_out = {8'd57, 8'd20, 1'b1, 1'b0};
119: data_out = {8'd58, 8'd20, 1'b1, 1'b0};
120: data_out = {8'd75, 8'd20, 1'b1, 1'b0};
121: data_out = {8'd76, 8'd20, 1'b1, 1'b0};
122: data_out = {8'd77, 8'd20, 1'b1, 1'b0};
123: data_out = {8'd78, 8'd20, 1'b1, 1'b0};
124: data_out = {8'd79, 8'd20, 1'b1, 1'b0};
125: data_out = {8'd80, 8'd20, 1'b1, 1'b0};
126: data_out = {8'd81, 8'd20, 1'b1, 1'b0};
127: data_out = {8'd82, 8'd20, 1'b1, 1'b0};
128: data_out = {8'd83, 8'd20, 1'b1, 1'b0};
129: data_out = {8'd84, 8'd20, 1'b1, 1'b0};
130: data_out = {8'd85, 8'd20, 1'b1, 1'b0};
131: data_out = {8'd86, 8'd20, 1'b1, 1'b0};
132: data_out = {8'd87, 8'd20, 1'b1, 1'b0};
133: data_out = {8'd88, 8'd20, 1'b1, 1'b0};
134: data_out = {8'd99, 8'd20, 1'b1, 1'b0};
135: data_out = {8'd100, 8'd20, 1'b1, 1'b0};
136: data_out = {8'd101, 8'd20, 1'b1, 1'b0};
137: data_out = {8'd102, 8'd20, 1'b1, 1'b0};
138: data_out = {8'd103, 8'd20, 1'b1, 1'b0};
139: data_out = {8'd104, 8'd20, 1'b1, 1'b0};
140: data_out = {8'd105, 8'd20, 1'b1, 1'b0};
141: data_out = {8'd106, 8'd20, 1'b1, 1'b0};
142: data_out = {8'd107, 8'd20, 1'b1, 1'b0};
143: data_out = {8'd108, 8'd20, 1'b1, 1'b0};
144: data_out = {8'd109, 8'd20, 1'b1, 1'b0};
145: data_out = {8'd110, 8'd20, 1'b1, 1'b0};
146: data_out = {8'd111, 8'd20, 1'b1, 1'b0};
147: data_out = {8'd112, 8'd20, 1'b1, 1'b0};
148: data_out = {8'd113, 8'd20, 1'b1, 1'b0};
149: data_out = {8'd114, 8'd20, 1'b1, 1'b0};
150: data_out = {8'd115, 8'd20, 1'b1, 1'b0};
151: data_out = {8'd116, 8'd20, 1'b1, 1'b0};
152: data_out = {8'd117, 8'd20, 1'b1, 1'b0};
153: data_out = {8'd118, 8'd20, 1'b1, 1'b0};
154: data_out = {8'd119, 8'd20, 1'b1, 1'b0};
155: data_out = {8'd129, 8'd20, 1'b1, 1'b0};
156: data_out = {8'd130, 8'd20, 1'b1, 1'b0};
157: data_out = {8'd131, 8'd20, 1'b1, 1'b0};
158: data_out = {8'd132, 8'd20, 1'b1, 1'b0};
159: data_out = {8'd133, 8'd20, 1'b1, 1'b0};
160: data_out = {8'd134, 8'd20, 1'b1, 1'b0};
161: data_out = {8'd135, 8'd20, 1'b1, 1'b0};
162: data_out = {8'd136, 8'd20, 1'b1, 1'b0};
163: data_out = {8'd137, 8'd20, 1'b1, 1'b0};
164: data_out = {8'd138, 8'd20, 1'b1, 1'b0};
165: data_out = {8'd139, 8'd20, 1'b1, 1'b0};
166: data_out = {8'd140, 8'd20, 1'b1, 1'b0};
167: data_out = {8'd141, 8'd20, 1'b1, 1'b0};
168: data_out = {8'd142, 8'd20, 1'b1, 1'b0};
169: data_out = {8'd143, 8'd20, 1'b1, 1'b0};
170: data_out = {8'd144, 8'd20, 1'b1, 1'b0};
171: data_out = {8'd145, 8'd20, 1'b1, 1'b0};
172: data_out = {8'd146, 8'd20, 1'b1, 1'b0};
173: data_out = {8'd147, 8'd20, 1'b1, 1'b0};
174: data_out = {8'd148, 8'd20, 1'b1, 1'b0};
175: data_out = {8'd149, 8'd20, 1'b1, 1'b0};
176: data_out = {8'd150, 8'd20, 1'b1, 1'b0};
177: data_out = {8'd151, 8'd20, 1'b1, 1'b0};
178: data_out = {8'd189, 8'd20, 1'b1, 1'b0};
179: data_out = {8'd190, 8'd20, 1'b1, 1'b0};
180: data_out = {8'd191, 8'd20, 1'b1, 1'b0};
181: data_out = {8'd192, 8'd20, 1'b1, 1'b0};
182: data_out = {8'd193, 8'd20, 1'b1, 1'b0};
183: data_out = {8'd194, 8'd20, 1'b1, 1'b0};
184: data_out = {8'd195, 8'd20, 1'b1, 1'b0};
185: data_out = {8'd196, 8'd20, 1'b1, 1'b0};
186: data_out = {8'd197, 8'd20, 1'b1, 1'b0};
187: data_out = {8'd198, 8'd20, 1'b1, 1'b0};
188: data_out = {8'd199, 8'd20, 1'b1, 1'b0};
189: data_out = {8'd200, 8'd20, 1'b1, 1'b0};
190: data_out = {8'd201, 8'd20, 1'b1, 1'b0};
191: data_out = {8'd202, 8'd20, 1'b1, 1'b0};
192: data_out = {8'd203, 8'd20, 1'b1, 1'b0};
193: data_out = {8'd204, 8'd20, 1'b1, 1'b0};
194: data_out = {8'd205, 8'd20, 1'b1, 1'b0};
195: data_out = {8'd206, 8'd20, 1'b1, 1'b0};
196: data_out = {8'd207, 8'd20, 1'b1, 1'b0};
197: data_out = {8'd208, 8'd20, 1'b1, 1'b0};
198: data_out = {8'd209, 8'd20, 1'b1, 1'b0};
199: data_out = {8'd7, 8'd21, 1'b1, 1'b0};
200: data_out = {8'd8, 8'd21, 1'b1, 1'b0};
201: data_out = {8'd9, 8'd21, 1'b1, 1'b0};
202: data_out = {8'd10, 8'd21, 1'b1, 1'b0};
203: data_out = {8'd11, 8'd21, 1'b1, 1'b0};
204: data_out = {8'd12, 8'd21, 1'b1, 1'b0};
205: data_out = {8'd13, 8'd21, 1'b1, 1'b0};
206: data_out = {8'd14, 8'd21, 1'b1, 1'b0};
207: data_out = {8'd15, 8'd21, 1'b1, 1'b0};
208: data_out = {8'd16, 8'd21, 1'b1, 1'b0};
209: data_out = {8'd17, 8'd21, 1'b1, 1'b0};
210: data_out = {8'd18, 8'd21, 1'b1, 1'b0};
211: data_out = {8'd19, 8'd21, 1'b1, 1'b0};
212: data_out = {8'd20, 8'd21, 1'b1, 1'b0};
213: data_out = {8'd21, 8'd21, 1'b1, 1'b0};
214: data_out = {8'd22, 8'd21, 1'b1, 1'b0};
215: data_out = {8'd23, 8'd21, 1'b1, 1'b0};
216: data_out = {8'd24, 8'd21, 1'b1, 1'b0};
217: data_out = {8'd25, 8'd21, 1'b1, 1'b0};
218: data_out = {8'd26, 8'd21, 1'b1, 1'b0};
219: data_out = {8'd27, 8'd21, 1'b1, 1'b0};
220: data_out = {8'd28, 8'd21, 1'b1, 1'b0};
221: data_out = {8'd29, 8'd21, 1'b1, 1'b0};
222: data_out = {8'd37, 8'd21, 1'b1, 1'b0};
223: data_out = {8'd38, 8'd21, 1'b1, 1'b0};
224: data_out = {8'd39, 8'd21, 1'b1, 1'b0};
225: data_out = {8'd40, 8'd21, 1'b1, 1'b0};
226: data_out = {8'd41, 8'd21, 1'b1, 1'b0};
227: data_out = {8'd42, 8'd21, 1'b1, 1'b0};
228: data_out = {8'd43, 8'd21, 1'b1, 1'b0};
229: data_out = {8'd44, 8'd21, 1'b1, 1'b0};
230: data_out = {8'd45, 8'd21, 1'b1, 1'b0};
231: data_out = {8'd46, 8'd21, 1'b1, 1'b0};
232: data_out = {8'd47, 8'd21, 1'b1, 1'b0};
233: data_out = {8'd48, 8'd21, 1'b1, 1'b0};
234: data_out = {8'd49, 8'd21, 1'b1, 1'b0};
235: data_out = {8'd50, 8'd21, 1'b1, 1'b0};
236: data_out = {8'd51, 8'd21, 1'b1, 1'b0};
237: data_out = {8'd52, 8'd21, 1'b1, 1'b0};
238: data_out = {8'd53, 8'd21, 1'b1, 1'b0};
239: data_out = {8'd54, 8'd21, 1'b1, 1'b0};
240: data_out = {8'd55, 8'd21, 1'b1, 1'b0};
241: data_out = {8'd56, 8'd21, 1'b1, 1'b0};
242: data_out = {8'd57, 8'd21, 1'b1, 1'b0};
243: data_out = {8'd58, 8'd21, 1'b1, 1'b0};
244: data_out = {8'd59, 8'd21, 1'b1, 1'b0};
245: data_out = {8'd74, 8'd21, 1'b1, 1'b0};
246: data_out = {8'd75, 8'd21, 1'b1, 1'b0};
247: data_out = {8'd76, 8'd21, 1'b1, 1'b0};
248: data_out = {8'd77, 8'd21, 1'b1, 1'b0};
249: data_out = {8'd78, 8'd21, 1'b1, 1'b0};
250: data_out = {8'd79, 8'd21, 1'b1, 1'b0};
251: data_out = {8'd80, 8'd21, 1'b1, 1'b0};
252: data_out = {8'd81, 8'd21, 1'b1, 1'b0};
253: data_out = {8'd82, 8'd21, 1'b1, 1'b0};
254: data_out = {8'd83, 8'd21, 1'b1, 1'b0};
255: data_out = {8'd84, 8'd21, 1'b1, 1'b0};
256: data_out = {8'd85, 8'd21, 1'b1, 1'b0};
257: data_out = {8'd86, 8'd21, 1'b1, 1'b0};
258: data_out = {8'd87, 8'd21, 1'b1, 1'b0};
259: data_out = {8'd88, 8'd21, 1'b1, 1'b0};
260: data_out = {8'd89, 8'd21, 1'b1, 1'b0};
261: data_out = {8'd98, 8'd21, 1'b1, 1'b0};
262: data_out = {8'd99, 8'd21, 1'b1, 1'b0};
263: data_out = {8'd100, 8'd21, 1'b1, 1'b0};
264: data_out = {8'd101, 8'd21, 1'b1, 1'b0};
265: data_out = {8'd102, 8'd21, 1'b1, 1'b0};
266: data_out = {8'd103, 8'd21, 1'b1, 1'b0};
267: data_out = {8'd104, 8'd21, 1'b1, 1'b0};
268: data_out = {8'd105, 8'd21, 1'b1, 1'b0};
269: data_out = {8'd106, 8'd21, 1'b1, 1'b0};
270: data_out = {8'd107, 8'd21, 1'b1, 1'b0};
271: data_out = {8'd108, 8'd21, 1'b1, 1'b0};
272: data_out = {8'd109, 8'd21, 1'b1, 1'b0};
273: data_out = {8'd110, 8'd21, 1'b1, 1'b0};
274: data_out = {8'd111, 8'd21, 1'b1, 1'b0};
275: data_out = {8'd112, 8'd21, 1'b1, 1'b0};
276: data_out = {8'd113, 8'd21, 1'b1, 1'b0};
277: data_out = {8'd114, 8'd21, 1'b1, 1'b0};
278: data_out = {8'd115, 8'd21, 1'b1, 1'b0};
279: data_out = {8'd116, 8'd21, 1'b1, 1'b0};
280: data_out = {8'd117, 8'd21, 1'b1, 1'b0};
281: data_out = {8'd118, 8'd21, 1'b1, 1'b0};
282: data_out = {8'd119, 8'd21, 1'b1, 1'b0};
283: data_out = {8'd120, 8'd21, 1'b1, 1'b0};
284: data_out = {8'd128, 8'd21, 1'b1, 1'b0};
285: data_out = {8'd129, 8'd21, 1'b1, 1'b0};
286: data_out = {8'd130, 8'd21, 1'b1, 1'b0};
287: data_out = {8'd131, 8'd21, 1'b1, 1'b0};
288: data_out = {8'd132, 8'd21, 1'b1, 1'b0};
289: data_out = {8'd133, 8'd21, 1'b1, 1'b0};
290: data_out = {8'd134, 8'd21, 1'b1, 1'b0};
291: data_out = {8'd135, 8'd21, 1'b1, 1'b0};
292: data_out = {8'd136, 8'd21, 1'b1, 1'b0};
293: data_out = {8'd137, 8'd21, 1'b1, 1'b0};
294: data_out = {8'd138, 8'd21, 1'b1, 1'b0};
295: data_out = {8'd139, 8'd21, 1'b1, 1'b0};
296: data_out = {8'd140, 8'd21, 1'b1, 1'b0};
297: data_out = {8'd141, 8'd21, 1'b1, 1'b0};
298: data_out = {8'd142, 8'd21, 1'b1, 1'b0};
299: data_out = {8'd143, 8'd21, 1'b1, 1'b0};
300: data_out = {8'd144, 8'd21, 1'b1, 1'b0};
301: data_out = {8'd145, 8'd21, 1'b1, 1'b0};
302: data_out = {8'd146, 8'd21, 1'b1, 1'b0};
303: data_out = {8'd147, 8'd21, 1'b1, 1'b0};
304: data_out = {8'd148, 8'd21, 1'b1, 1'b0};
305: data_out = {8'd149, 8'd21, 1'b1, 1'b0};
306: data_out = {8'd150, 8'd21, 1'b1, 1'b0};
307: data_out = {8'd151, 8'd21, 1'b1, 1'b0};
308: data_out = {8'd188, 8'd21, 1'b1, 1'b0};
309: data_out = {8'd189, 8'd21, 1'b1, 1'b0};
310: data_out = {8'd190, 8'd21, 1'b1, 1'b0};
311: data_out = {8'd191, 8'd21, 1'b1, 1'b0};
312: data_out = {8'd192, 8'd21, 1'b1, 1'b0};
313: data_out = {8'd193, 8'd21, 1'b1, 1'b0};
314: data_out = {8'd194, 8'd21, 1'b1, 1'b0};
315: data_out = {8'd195, 8'd21, 1'b1, 1'b0};
316: data_out = {8'd196, 8'd21, 1'b1, 1'b0};
317: data_out = {8'd197, 8'd21, 1'b1, 1'b0};
318: data_out = {8'd198, 8'd21, 1'b1, 1'b0};
319: data_out = {8'd199, 8'd21, 1'b1, 1'b0};
320: data_out = {8'd200, 8'd21, 1'b1, 1'b0};
321: data_out = {8'd201, 8'd21, 1'b1, 1'b0};
322: data_out = {8'd202, 8'd21, 1'b1, 1'b0};
323: data_out = {8'd203, 8'd21, 1'b1, 1'b0};
324: data_out = {8'd204, 8'd21, 1'b1, 1'b0};
325: data_out = {8'd205, 8'd21, 1'b1, 1'b0};
326: data_out = {8'd206, 8'd21, 1'b1, 1'b0};
327: data_out = {8'd207, 8'd21, 1'b1, 1'b0};
328: data_out = {8'd208, 8'd21, 1'b1, 1'b0};
329: data_out = {8'd209, 8'd21, 1'b1, 1'b0};
330: data_out = {8'd210, 8'd21, 1'b1, 1'b0};
331: data_out = {8'd6, 8'd22, 1'b1, 1'b0};
332: data_out = {8'd7, 8'd22, 1'b1, 1'b0};
333: data_out = {8'd8, 8'd22, 1'b1, 1'b0};
334: data_out = {8'd9, 8'd22, 1'b1, 1'b0};
335: data_out = {8'd10, 8'd22, 1'b1, 1'b0};
336: data_out = {8'd11, 8'd22, 1'b1, 1'b0};
337: data_out = {8'd12, 8'd22, 1'b1, 1'b0};
338: data_out = {8'd13, 8'd22, 1'b1, 1'b0};
339: data_out = {8'd14, 8'd22, 1'b1, 1'b0};
340: data_out = {8'd15, 8'd22, 1'b1, 1'b0};
341: data_out = {8'd16, 8'd22, 1'b1, 1'b0};
342: data_out = {8'd17, 8'd22, 1'b1, 1'b0};
343: data_out = {8'd18, 8'd22, 1'b1, 1'b0};
344: data_out = {8'd19, 8'd22, 1'b1, 1'b0};
345: data_out = {8'd20, 8'd22, 1'b1, 1'b0};
346: data_out = {8'd21, 8'd22, 1'b1, 1'b0};
347: data_out = {8'd22, 8'd22, 1'b1, 1'b0};
348: data_out = {8'd23, 8'd22, 1'b1, 1'b0};
349: data_out = {8'd24, 8'd22, 1'b1, 1'b0};
350: data_out = {8'd25, 8'd22, 1'b1, 1'b0};
351: data_out = {8'd26, 8'd22, 1'b1, 1'b0};
352: data_out = {8'd27, 8'd22, 1'b1, 1'b0};
353: data_out = {8'd28, 8'd22, 1'b1, 1'b0};
354: data_out = {8'd29, 8'd22, 1'b1, 1'b0};
355: data_out = {8'd30, 8'd22, 1'b1, 1'b0};
356: data_out = {8'd36, 8'd22, 1'b1, 1'b0};
357: data_out = {8'd37, 8'd22, 1'b1, 1'b0};
358: data_out = {8'd38, 8'd22, 1'b1, 1'b0};
359: data_out = {8'd39, 8'd22, 1'b1, 1'b0};
360: data_out = {8'd40, 8'd22, 1'b1, 1'b0};
361: data_out = {8'd41, 8'd22, 1'b1, 1'b0};
362: data_out = {8'd42, 8'd22, 1'b1, 1'b0};
363: data_out = {8'd43, 8'd22, 1'b1, 1'b0};
364: data_out = {8'd44, 8'd22, 1'b1, 1'b0};
365: data_out = {8'd45, 8'd22, 1'b1, 1'b0};
366: data_out = {8'd46, 8'd22, 1'b1, 1'b0};
367: data_out = {8'd47, 8'd22, 1'b1, 1'b0};
368: data_out = {8'd48, 8'd22, 1'b1, 1'b0};
369: data_out = {8'd49, 8'd22, 1'b1, 1'b0};
370: data_out = {8'd50, 8'd22, 1'b1, 1'b0};
371: data_out = {8'd51, 8'd22, 1'b1, 1'b0};
372: data_out = {8'd52, 8'd22, 1'b1, 1'b0};
373: data_out = {8'd53, 8'd22, 1'b1, 1'b0};
374: data_out = {8'd54, 8'd22, 1'b1, 1'b0};
375: data_out = {8'd55, 8'd22, 1'b1, 1'b0};
376: data_out = {8'd56, 8'd22, 1'b1, 1'b0};
377: data_out = {8'd57, 8'd22, 1'b1, 1'b0};
378: data_out = {8'd58, 8'd22, 1'b1, 1'b0};
379: data_out = {8'd59, 8'd22, 1'b1, 1'b0};
380: data_out = {8'd60, 8'd22, 1'b1, 1'b0};
381: data_out = {8'd73, 8'd22, 1'b1, 1'b0};
382: data_out = {8'd74, 8'd22, 1'b1, 1'b0};
383: data_out = {8'd75, 8'd22, 1'b1, 1'b0};
384: data_out = {8'd76, 8'd22, 1'b1, 1'b0};
385: data_out = {8'd77, 8'd22, 1'b1, 1'b0};
386: data_out = {8'd78, 8'd22, 1'b1, 1'b0};
387: data_out = {8'd79, 8'd22, 1'b1, 1'b0};
388: data_out = {8'd80, 8'd22, 1'b1, 1'b0};
389: data_out = {8'd81, 8'd22, 1'b1, 1'b0};
390: data_out = {8'd82, 8'd22, 1'b1, 1'b0};
391: data_out = {8'd83, 8'd22, 1'b1, 1'b0};
392: data_out = {8'd84, 8'd22, 1'b1, 1'b0};
393: data_out = {8'd85, 8'd22, 1'b1, 1'b0};
394: data_out = {8'd86, 8'd22, 1'b1, 1'b0};
395: data_out = {8'd87, 8'd22, 1'b1, 1'b0};
396: data_out = {8'd88, 8'd22, 1'b1, 1'b0};
397: data_out = {8'd89, 8'd22, 1'b1, 1'b0};
398: data_out = {8'd90, 8'd22, 1'b1, 1'b0};
399: data_out = {8'd97, 8'd22, 1'b1, 1'b0};
400: data_out = {8'd98, 8'd22, 1'b1, 1'b0};
401: data_out = {8'd99, 8'd22, 1'b1, 1'b0};
402: data_out = {8'd100, 8'd22, 1'b1, 1'b0};
403: data_out = {8'd101, 8'd22, 1'b1, 1'b0};
404: data_out = {8'd102, 8'd22, 1'b1, 1'b0};
405: data_out = {8'd103, 8'd22, 1'b1, 1'b0};
406: data_out = {8'd104, 8'd22, 1'b1, 1'b0};
407: data_out = {8'd105, 8'd22, 1'b1, 1'b0};
408: data_out = {8'd106, 8'd22, 1'b1, 1'b0};
409: data_out = {8'd107, 8'd22, 1'b1, 1'b0};
410: data_out = {8'd108, 8'd22, 1'b1, 1'b0};
411: data_out = {8'd109, 8'd22, 1'b1, 1'b0};
412: data_out = {8'd110, 8'd22, 1'b1, 1'b0};
413: data_out = {8'd111, 8'd22, 1'b1, 1'b0};
414: data_out = {8'd112, 8'd22, 1'b1, 1'b0};
415: data_out = {8'd113, 8'd22, 1'b1, 1'b0};
416: data_out = {8'd114, 8'd22, 1'b1, 1'b0};
417: data_out = {8'd115, 8'd22, 1'b1, 1'b0};
418: data_out = {8'd116, 8'd22, 1'b1, 1'b0};
419: data_out = {8'd117, 8'd22, 1'b1, 1'b0};
420: data_out = {8'd118, 8'd22, 1'b1, 1'b0};
421: data_out = {8'd119, 8'd22, 1'b1, 1'b0};
422: data_out = {8'd120, 8'd22, 1'b1, 1'b0};
423: data_out = {8'd121, 8'd22, 1'b1, 1'b0};
424: data_out = {8'd127, 8'd22, 1'b1, 1'b0};
425: data_out = {8'd128, 8'd22, 1'b1, 1'b0};
426: data_out = {8'd129, 8'd22, 1'b1, 1'b0};
427: data_out = {8'd130, 8'd22, 1'b1, 1'b0};
428: data_out = {8'd131, 8'd22, 1'b1, 1'b0};
429: data_out = {8'd132, 8'd22, 1'b1, 1'b0};
430: data_out = {8'd133, 8'd22, 1'b1, 1'b0};
431: data_out = {8'd134, 8'd22, 1'b1, 1'b0};
432: data_out = {8'd135, 8'd22, 1'b1, 1'b0};
433: data_out = {8'd136, 8'd22, 1'b1, 1'b0};
434: data_out = {8'd137, 8'd22, 1'b1, 1'b0};
435: data_out = {8'd138, 8'd22, 1'b1, 1'b0};
436: data_out = {8'd139, 8'd22, 1'b1, 1'b0};
437: data_out = {8'd140, 8'd22, 1'b1, 1'b0};
438: data_out = {8'd141, 8'd22, 1'b1, 1'b0};
439: data_out = {8'd142, 8'd22, 1'b1, 1'b0};
440: data_out = {8'd143, 8'd22, 1'b1, 1'b0};
441: data_out = {8'd144, 8'd22, 1'b1, 1'b0};
442: data_out = {8'd145, 8'd22, 1'b1, 1'b0};
443: data_out = {8'd146, 8'd22, 1'b1, 1'b0};
444: data_out = {8'd147, 8'd22, 1'b1, 1'b0};
445: data_out = {8'd148, 8'd22, 1'b1, 1'b0};
446: data_out = {8'd149, 8'd22, 1'b1, 1'b0};
447: data_out = {8'd150, 8'd22, 1'b1, 1'b0};
448: data_out = {8'd151, 8'd22, 1'b1, 1'b0};
449: data_out = {8'd187, 8'd22, 1'b1, 1'b0};
450: data_out = {8'd188, 8'd22, 1'b1, 1'b0};
451: data_out = {8'd189, 8'd22, 1'b1, 1'b0};
452: data_out = {8'd190, 8'd22, 1'b1, 1'b0};
453: data_out = {8'd191, 8'd22, 1'b1, 1'b0};
454: data_out = {8'd192, 8'd22, 1'b1, 1'b0};
455: data_out = {8'd193, 8'd22, 1'b1, 1'b0};
456: data_out = {8'd194, 8'd22, 1'b1, 1'b0};
457: data_out = {8'd195, 8'd22, 1'b1, 1'b0};
458: data_out = {8'd196, 8'd22, 1'b1, 1'b0};
459: data_out = {8'd197, 8'd22, 1'b1, 1'b0};
460: data_out = {8'd198, 8'd22, 1'b1, 1'b0};
461: data_out = {8'd199, 8'd22, 1'b1, 1'b0};
462: data_out = {8'd200, 8'd22, 1'b1, 1'b0};
463: data_out = {8'd201, 8'd22, 1'b1, 1'b0};
464: data_out = {8'd202, 8'd22, 1'b1, 1'b0};
465: data_out = {8'd203, 8'd22, 1'b1, 1'b0};
466: data_out = {8'd204, 8'd22, 1'b1, 1'b0};
467: data_out = {8'd205, 8'd22, 1'b1, 1'b0};
468: data_out = {8'd206, 8'd22, 1'b1, 1'b0};
469: data_out = {8'd207, 8'd22, 1'b1, 1'b0};
470: data_out = {8'd208, 8'd22, 1'b1, 1'b0};
471: data_out = {8'd209, 8'd22, 1'b1, 1'b0};
472: data_out = {8'd210, 8'd22, 1'b1, 1'b0};
473: data_out = {8'd211, 8'd22, 1'b1, 1'b0};
474: data_out = {8'd6, 8'd23, 1'b1, 1'b0};
475: data_out = {8'd7, 8'd23, 1'b1, 1'b0};
476: data_out = {8'd8, 8'd23, 1'b1, 1'b0};
477: data_out = {8'd9, 8'd23, 1'b1, 1'b0};
478: data_out = {8'd10, 8'd23, 1'b1, 1'b0};
479: data_out = {8'd11, 8'd23, 1'b1, 1'b0};
480: data_out = {8'd12, 8'd23, 1'b1, 1'b0};
481: data_out = {8'd13, 8'd23, 1'b1, 1'b0};
482: data_out = {8'd14, 8'd23, 1'b1, 1'b0};
483: data_out = {8'd15, 8'd23, 1'b1, 1'b0};
484: data_out = {8'd16, 8'd23, 1'b1, 1'b0};
485: data_out = {8'd17, 8'd23, 1'b1, 1'b0};
486: data_out = {8'd18, 8'd23, 1'b1, 1'b0};
487: data_out = {8'd19, 8'd23, 1'b1, 1'b0};
488: data_out = {8'd20, 8'd23, 1'b1, 1'b0};
489: data_out = {8'd21, 8'd23, 1'b1, 1'b0};
490: data_out = {8'd22, 8'd23, 1'b1, 1'b0};
491: data_out = {8'd23, 8'd23, 1'b1, 1'b0};
492: data_out = {8'd24, 8'd23, 1'b1, 1'b0};
493: data_out = {8'd25, 8'd23, 1'b1, 1'b0};
494: data_out = {8'd26, 8'd23, 1'b1, 1'b0};
495: data_out = {8'd27, 8'd23, 1'b1, 1'b0};
496: data_out = {8'd28, 8'd23, 1'b1, 1'b0};
497: data_out = {8'd29, 8'd23, 1'b1, 1'b0};
498: data_out = {8'd30, 8'd23, 1'b1, 1'b0};
499: data_out = {8'd36, 8'd23, 1'b1, 1'b0};
500: data_out = {8'd37, 8'd23, 1'b1, 1'b0};
501: data_out = {8'd38, 8'd23, 1'b1, 1'b0};
502: data_out = {8'd39, 8'd23, 1'b1, 1'b0};
503: data_out = {8'd40, 8'd23, 1'b1, 1'b0};
504: data_out = {8'd41, 8'd23, 1'b1, 1'b0};
505: data_out = {8'd42, 8'd23, 1'b1, 1'b0};
506: data_out = {8'd43, 8'd23, 1'b1, 1'b0};
507: data_out = {8'd44, 8'd23, 1'b1, 1'b0};
508: data_out = {8'd45, 8'd23, 1'b1, 1'b0};
509: data_out = {8'd46, 8'd23, 1'b1, 1'b0};
510: data_out = {8'd47, 8'd23, 1'b1, 1'b0};
511: data_out = {8'd48, 8'd23, 1'b1, 1'b0};
512: data_out = {8'd49, 8'd23, 1'b1, 1'b0};
513: data_out = {8'd50, 8'd23, 1'b1, 1'b0};
514: data_out = {8'd51, 8'd23, 1'b1, 1'b0};
515: data_out = {8'd52, 8'd23, 1'b1, 1'b0};
516: data_out = {8'd53, 8'd23, 1'b1, 1'b0};
517: data_out = {8'd54, 8'd23, 1'b1, 1'b0};
518: data_out = {8'd55, 8'd23, 1'b1, 1'b0};
519: data_out = {8'd56, 8'd23, 1'b1, 1'b0};
520: data_out = {8'd57, 8'd23, 1'b1, 1'b0};
521: data_out = {8'd58, 8'd23, 1'b1, 1'b0};
522: data_out = {8'd59, 8'd23, 1'b1, 1'b0};
523: data_out = {8'd60, 8'd23, 1'b1, 1'b0};
524: data_out = {8'd73, 8'd23, 1'b1, 1'b0};
525: data_out = {8'd74, 8'd23, 1'b1, 1'b0};
526: data_out = {8'd75, 8'd23, 1'b1, 1'b0};
527: data_out = {8'd76, 8'd23, 1'b1, 1'b0};
528: data_out = {8'd77, 8'd23, 1'b1, 1'b0};
529: data_out = {8'd78, 8'd23, 1'b1, 1'b0};
530: data_out = {8'd79, 8'd23, 1'b1, 1'b0};
531: data_out = {8'd80, 8'd23, 1'b1, 1'b0};
532: data_out = {8'd81, 8'd23, 1'b1, 1'b0};
533: data_out = {8'd82, 8'd23, 1'b1, 1'b0};
534: data_out = {8'd83, 8'd23, 1'b1, 1'b0};
535: data_out = {8'd84, 8'd23, 1'b1, 1'b0};
536: data_out = {8'd85, 8'd23, 1'b1, 1'b0};
537: data_out = {8'd86, 8'd23, 1'b1, 1'b0};
538: data_out = {8'd87, 8'd23, 1'b1, 1'b0};
539: data_out = {8'd88, 8'd23, 1'b1, 1'b0};
540: data_out = {8'd89, 8'd23, 1'b1, 1'b0};
541: data_out = {8'd90, 8'd23, 1'b1, 1'b0};
542: data_out = {8'd97, 8'd23, 1'b1, 1'b0};
543: data_out = {8'd98, 8'd23, 1'b1, 1'b0};
544: data_out = {8'd99, 8'd23, 1'b1, 1'b0};
545: data_out = {8'd100, 8'd23, 1'b1, 1'b0};
546: data_out = {8'd101, 8'd23, 1'b1, 1'b0};
547: data_out = {8'd102, 8'd23, 1'b1, 1'b0};
548: data_out = {8'd103, 8'd23, 1'b1, 1'b0};
549: data_out = {8'd104, 8'd23, 1'b1, 1'b0};
550: data_out = {8'd105, 8'd23, 1'b1, 1'b0};
551: data_out = {8'd106, 8'd23, 1'b1, 1'b0};
552: data_out = {8'd107, 8'd23, 1'b1, 1'b0};
553: data_out = {8'd108, 8'd23, 1'b1, 1'b0};
554: data_out = {8'd109, 8'd23, 1'b1, 1'b0};
555: data_out = {8'd110, 8'd23, 1'b1, 1'b0};
556: data_out = {8'd111, 8'd23, 1'b1, 1'b0};
557: data_out = {8'd112, 8'd23, 1'b1, 1'b0};
558: data_out = {8'd113, 8'd23, 1'b1, 1'b0};
559: data_out = {8'd114, 8'd23, 1'b1, 1'b0};
560: data_out = {8'd115, 8'd23, 1'b1, 1'b0};
561: data_out = {8'd116, 8'd23, 1'b1, 1'b0};
562: data_out = {8'd117, 8'd23, 1'b1, 1'b0};
563: data_out = {8'd118, 8'd23, 1'b1, 1'b0};
564: data_out = {8'd119, 8'd23, 1'b1, 1'b0};
565: data_out = {8'd120, 8'd23, 1'b1, 1'b0};
566: data_out = {8'd121, 8'd23, 1'b1, 1'b0};
567: data_out = {8'd127, 8'd23, 1'b1, 1'b0};
568: data_out = {8'd128, 8'd23, 1'b1, 1'b0};
569: data_out = {8'd129, 8'd23, 1'b1, 1'b0};
570: data_out = {8'd130, 8'd23, 1'b1, 1'b0};
571: data_out = {8'd131, 8'd23, 1'b1, 1'b0};
572: data_out = {8'd132, 8'd23, 1'b1, 1'b0};
573: data_out = {8'd133, 8'd23, 1'b1, 1'b0};
574: data_out = {8'd134, 8'd23, 1'b1, 1'b0};
575: data_out = {8'd135, 8'd23, 1'b1, 1'b0};
576: data_out = {8'd136, 8'd23, 1'b1, 1'b0};
577: data_out = {8'd137, 8'd23, 1'b1, 1'b0};
578: data_out = {8'd138, 8'd23, 1'b1, 1'b0};
579: data_out = {8'd139, 8'd23, 1'b1, 1'b0};
580: data_out = {8'd140, 8'd23, 1'b1, 1'b0};
581: data_out = {8'd141, 8'd23, 1'b1, 1'b0};
582: data_out = {8'd142, 8'd23, 1'b1, 1'b0};
583: data_out = {8'd143, 8'd23, 1'b1, 1'b0};
584: data_out = {8'd144, 8'd23, 1'b1, 1'b0};
585: data_out = {8'd145, 8'd23, 1'b1, 1'b0};
586: data_out = {8'd146, 8'd23, 1'b1, 1'b0};
587: data_out = {8'd147, 8'd23, 1'b1, 1'b0};
588: data_out = {8'd148, 8'd23, 1'b1, 1'b0};
589: data_out = {8'd149, 8'd23, 1'b1, 1'b0};
590: data_out = {8'd150, 8'd23, 1'b1, 1'b0};
591: data_out = {8'd151, 8'd23, 1'b1, 1'b0};
592: data_out = {8'd187, 8'd23, 1'b1, 1'b0};
593: data_out = {8'd188, 8'd23, 1'b1, 1'b0};
594: data_out = {8'd189, 8'd23, 1'b1, 1'b0};
595: data_out = {8'd190, 8'd23, 1'b1, 1'b0};
596: data_out = {8'd191, 8'd23, 1'b1, 1'b0};
597: data_out = {8'd192, 8'd23, 1'b1, 1'b0};
598: data_out = {8'd193, 8'd23, 1'b1, 1'b0};
599: data_out = {8'd194, 8'd23, 1'b1, 1'b0};
600: data_out = {8'd195, 8'd23, 1'b1, 1'b0};
601: data_out = {8'd196, 8'd23, 1'b1, 1'b0};
602: data_out = {8'd197, 8'd23, 1'b1, 1'b0};
603: data_out = {8'd198, 8'd23, 1'b1, 1'b0};
604: data_out = {8'd199, 8'd23, 1'b1, 1'b0};
605: data_out = {8'd200, 8'd23, 1'b1, 1'b0};
606: data_out = {8'd201, 8'd23, 1'b1, 1'b0};
607: data_out = {8'd202, 8'd23, 1'b1, 1'b0};
608: data_out = {8'd203, 8'd23, 1'b1, 1'b0};
609: data_out = {8'd204, 8'd23, 1'b1, 1'b0};
610: data_out = {8'd205, 8'd23, 1'b1, 1'b0};
611: data_out = {8'd206, 8'd23, 1'b1, 1'b0};
612: data_out = {8'd207, 8'd23, 1'b1, 1'b0};
613: data_out = {8'd208, 8'd23, 1'b1, 1'b0};
614: data_out = {8'd209, 8'd23, 1'b1, 1'b0};
615: data_out = {8'd210, 8'd23, 1'b1, 1'b0};
616: data_out = {8'd211, 8'd23, 1'b1, 1'b0};
617: data_out = {8'd6, 8'd24, 1'b1, 1'b0};
618: data_out = {8'd7, 8'd24, 1'b1, 1'b0};
619: data_out = {8'd8, 8'd24, 1'b1, 1'b0};
620: data_out = {8'd9, 8'd24, 1'b1, 1'b0};
621: data_out = {8'd10, 8'd24, 1'b1, 1'b0};
622: data_out = {8'd11, 8'd24, 1'b1, 1'b0};
623: data_out = {8'd12, 8'd24, 1'b1, 1'b0};
624: data_out = {8'd13, 8'd24, 1'b1, 1'b0};
625: data_out = {8'd14, 8'd24, 1'b1, 1'b0};
626: data_out = {8'd15, 8'd24, 1'b1, 1'b0};
627: data_out = {8'd16, 8'd24, 1'b1, 1'b0};
628: data_out = {8'd17, 8'd24, 1'b1, 1'b0};
629: data_out = {8'd18, 8'd24, 1'b1, 1'b0};
630: data_out = {8'd19, 8'd24, 1'b1, 1'b0};
631: data_out = {8'd20, 8'd24, 1'b1, 1'b0};
632: data_out = {8'd21, 8'd24, 1'b1, 1'b0};
633: data_out = {8'd22, 8'd24, 1'b1, 1'b0};
634: data_out = {8'd23, 8'd24, 1'b1, 1'b0};
635: data_out = {8'd24, 8'd24, 1'b1, 1'b0};
636: data_out = {8'd25, 8'd24, 1'b1, 1'b0};
637: data_out = {8'd26, 8'd24, 1'b1, 1'b0};
638: data_out = {8'd27, 8'd24, 1'b1, 1'b0};
639: data_out = {8'd28, 8'd24, 1'b1, 1'b0};
640: data_out = {8'd29, 8'd24, 1'b1, 1'b0};
641: data_out = {8'd30, 8'd24, 1'b1, 1'b0};
642: data_out = {8'd36, 8'd24, 1'b1, 1'b0};
643: data_out = {8'd37, 8'd24, 1'b1, 1'b0};
644: data_out = {8'd38, 8'd24, 1'b1, 1'b0};
645: data_out = {8'd39, 8'd24, 1'b1, 1'b0};
646: data_out = {8'd40, 8'd24, 1'b1, 1'b0};
647: data_out = {8'd41, 8'd24, 1'b1, 1'b0};
648: data_out = {8'd42, 8'd24, 1'b1, 1'b0};
649: data_out = {8'd43, 8'd24, 1'b1, 1'b0};
650: data_out = {8'd44, 8'd24, 1'b1, 1'b0};
651: data_out = {8'd45, 8'd24, 1'b1, 1'b0};
652: data_out = {8'd46, 8'd24, 1'b1, 1'b0};
653: data_out = {8'd47, 8'd24, 1'b1, 1'b0};
654: data_out = {8'd48, 8'd24, 1'b1, 1'b0};
655: data_out = {8'd49, 8'd24, 1'b1, 1'b0};
656: data_out = {8'd50, 8'd24, 1'b1, 1'b0};
657: data_out = {8'd51, 8'd24, 1'b1, 1'b0};
658: data_out = {8'd52, 8'd24, 1'b1, 1'b0};
659: data_out = {8'd53, 8'd24, 1'b1, 1'b0};
660: data_out = {8'd54, 8'd24, 1'b1, 1'b0};
661: data_out = {8'd55, 8'd24, 1'b1, 1'b0};
662: data_out = {8'd56, 8'd24, 1'b1, 1'b0};
663: data_out = {8'd57, 8'd24, 1'b1, 1'b0};
664: data_out = {8'd58, 8'd24, 1'b1, 1'b0};
665: data_out = {8'd59, 8'd24, 1'b1, 1'b0};
666: data_out = {8'd60, 8'd24, 1'b1, 1'b0};
667: data_out = {8'd73, 8'd24, 1'b1, 1'b0};
668: data_out = {8'd74, 8'd24, 1'b1, 1'b0};
669: data_out = {8'd75, 8'd24, 1'b1, 1'b0};
670: data_out = {8'd76, 8'd24, 1'b1, 1'b0};
671: data_out = {8'd77, 8'd24, 1'b1, 1'b0};
672: data_out = {8'd78, 8'd24, 1'b1, 1'b0};
673: data_out = {8'd79, 8'd24, 1'b1, 1'b0};
674: data_out = {8'd80, 8'd24, 1'b1, 1'b0};
675: data_out = {8'd81, 8'd24, 1'b1, 1'b0};
676: data_out = {8'd82, 8'd24, 1'b1, 1'b0};
677: data_out = {8'd83, 8'd24, 1'b1, 1'b0};
678: data_out = {8'd84, 8'd24, 1'b1, 1'b0};
679: data_out = {8'd85, 8'd24, 1'b1, 1'b0};
680: data_out = {8'd86, 8'd24, 1'b1, 1'b0};
681: data_out = {8'd87, 8'd24, 1'b1, 1'b0};
682: data_out = {8'd88, 8'd24, 1'b1, 1'b0};
683: data_out = {8'd89, 8'd24, 1'b1, 1'b0};
684: data_out = {8'd90, 8'd24, 1'b1, 1'b0};
685: data_out = {8'd97, 8'd24, 1'b1, 1'b0};
686: data_out = {8'd98, 8'd24, 1'b1, 1'b0};
687: data_out = {8'd99, 8'd24, 1'b1, 1'b0};
688: data_out = {8'd100, 8'd24, 1'b1, 1'b0};
689: data_out = {8'd101, 8'd24, 1'b1, 1'b0};
690: data_out = {8'd102, 8'd24, 1'b1, 1'b0};
691: data_out = {8'd103, 8'd24, 1'b1, 1'b0};
692: data_out = {8'd104, 8'd24, 1'b1, 1'b0};
693: data_out = {8'd105, 8'd24, 1'b1, 1'b0};
694: data_out = {8'd106, 8'd24, 1'b1, 1'b0};
695: data_out = {8'd107, 8'd24, 1'b1, 1'b0};
696: data_out = {8'd108, 8'd24, 1'b1, 1'b0};
697: data_out = {8'd109, 8'd24, 1'b1, 1'b0};
698: data_out = {8'd110, 8'd24, 1'b1, 1'b0};
699: data_out = {8'd111, 8'd24, 1'b1, 1'b0};
700: data_out = {8'd112, 8'd24, 1'b1, 1'b0};
701: data_out = {8'd113, 8'd24, 1'b1, 1'b0};
702: data_out = {8'd114, 8'd24, 1'b1, 1'b0};
703: data_out = {8'd115, 8'd24, 1'b1, 1'b0};
704: data_out = {8'd116, 8'd24, 1'b1, 1'b0};
705: data_out = {8'd117, 8'd24, 1'b1, 1'b0};
706: data_out = {8'd118, 8'd24, 1'b1, 1'b0};
707: data_out = {8'd119, 8'd24, 1'b1, 1'b0};
708: data_out = {8'd120, 8'd24, 1'b1, 1'b0};
709: data_out = {8'd121, 8'd24, 1'b1, 1'b0};
710: data_out = {8'd127, 8'd24, 1'b1, 1'b0};
711: data_out = {8'd128, 8'd24, 1'b1, 1'b0};
712: data_out = {8'd129, 8'd24, 1'b1, 1'b0};
713: data_out = {8'd130, 8'd24, 1'b1, 1'b0};
714: data_out = {8'd131, 8'd24, 1'b1, 1'b0};
715: data_out = {8'd132, 8'd24, 1'b1, 1'b0};
716: data_out = {8'd133, 8'd24, 1'b1, 1'b0};
717: data_out = {8'd134, 8'd24, 1'b1, 1'b0};
718: data_out = {8'd135, 8'd24, 1'b1, 1'b0};
719: data_out = {8'd136, 8'd24, 1'b1, 1'b0};
720: data_out = {8'd137, 8'd24, 1'b1, 1'b0};
721: data_out = {8'd138, 8'd24, 1'b1, 1'b0};
722: data_out = {8'd139, 8'd24, 1'b1, 1'b0};
723: data_out = {8'd140, 8'd24, 1'b1, 1'b0};
724: data_out = {8'd141, 8'd24, 1'b1, 1'b0};
725: data_out = {8'd142, 8'd24, 1'b1, 1'b0};
726: data_out = {8'd143, 8'd24, 1'b1, 1'b0};
727: data_out = {8'd144, 8'd24, 1'b1, 1'b0};
728: data_out = {8'd145, 8'd24, 1'b1, 1'b0};
729: data_out = {8'd146, 8'd24, 1'b1, 1'b0};
730: data_out = {8'd147, 8'd24, 1'b1, 1'b0};
731: data_out = {8'd148, 8'd24, 1'b1, 1'b0};
732: data_out = {8'd149, 8'd24, 1'b1, 1'b0};
733: data_out = {8'd150, 8'd24, 1'b1, 1'b0};
734: data_out = {8'd151, 8'd24, 1'b1, 1'b0};
735: data_out = {8'd187, 8'd24, 1'b1, 1'b0};
736: data_out = {8'd188, 8'd24, 1'b1, 1'b0};
737: data_out = {8'd189, 8'd24, 1'b1, 1'b0};
738: data_out = {8'd190, 8'd24, 1'b1, 1'b0};
739: data_out = {8'd191, 8'd24, 1'b1, 1'b0};
740: data_out = {8'd192, 8'd24, 1'b1, 1'b0};
741: data_out = {8'd193, 8'd24, 1'b1, 1'b0};
742: data_out = {8'd194, 8'd24, 1'b1, 1'b0};
743: data_out = {8'd195, 8'd24, 1'b1, 1'b0};
744: data_out = {8'd196, 8'd24, 1'b1, 1'b0};
745: data_out = {8'd197, 8'd24, 1'b1, 1'b0};
746: data_out = {8'd198, 8'd24, 1'b1, 1'b0};
747: data_out = {8'd199, 8'd24, 1'b1, 1'b0};
748: data_out = {8'd200, 8'd24, 1'b1, 1'b0};
749: data_out = {8'd201, 8'd24, 1'b1, 1'b0};
750: data_out = {8'd202, 8'd24, 1'b1, 1'b0};
751: data_out = {8'd203, 8'd24, 1'b1, 1'b0};
752: data_out = {8'd204, 8'd24, 1'b1, 1'b0};
753: data_out = {8'd205, 8'd24, 1'b1, 1'b0};
754: data_out = {8'd206, 8'd24, 1'b1, 1'b0};
755: data_out = {8'd207, 8'd24, 1'b1, 1'b0};
756: data_out = {8'd208, 8'd24, 1'b1, 1'b0};
757: data_out = {8'd209, 8'd24, 1'b1, 1'b0};
758: data_out = {8'd210, 8'd24, 1'b1, 1'b0};
759: data_out = {8'd211, 8'd24, 1'b1, 1'b0};
760: data_out = {8'd6, 8'd25, 1'b1, 1'b0};
761: data_out = {8'd7, 8'd25, 1'b1, 1'b0};
762: data_out = {8'd8, 8'd25, 1'b1, 1'b0};
763: data_out = {8'd9, 8'd25, 1'b1, 1'b0};
764: data_out = {8'd10, 8'd25, 1'b1, 1'b0};
765: data_out = {8'd11, 8'd25, 1'b1, 1'b0};
766: data_out = {8'd25, 8'd25, 1'b1, 1'b0};
767: data_out = {8'd26, 8'd25, 1'b1, 1'b0};
768: data_out = {8'd27, 8'd25, 1'b1, 1'b0};
769: data_out = {8'd28, 8'd25, 1'b1, 1'b0};
770: data_out = {8'd29, 8'd25, 1'b1, 1'b0};
771: data_out = {8'd30, 8'd25, 1'b1, 1'b0};
772: data_out = {8'd36, 8'd25, 1'b1, 1'b0};
773: data_out = {8'd37, 8'd25, 1'b1, 1'b0};
774: data_out = {8'd38, 8'd25, 1'b1, 1'b0};
775: data_out = {8'd39, 8'd25, 1'b1, 1'b0};
776: data_out = {8'd40, 8'd25, 1'b1, 1'b0};
777: data_out = {8'd41, 8'd25, 1'b1, 1'b0};
778: data_out = {8'd55, 8'd25, 1'b1, 1'b0};
779: data_out = {8'd56, 8'd25, 1'b1, 1'b0};
780: data_out = {8'd57, 8'd25, 1'b1, 1'b0};
781: data_out = {8'd58, 8'd25, 1'b1, 1'b0};
782: data_out = {8'd59, 8'd25, 1'b1, 1'b0};
783: data_out = {8'd60, 8'd25, 1'b1, 1'b0};
784: data_out = {8'd73, 8'd25, 1'b1, 1'b0};
785: data_out = {8'd74, 8'd25, 1'b1, 1'b0};
786: data_out = {8'd75, 8'd25, 1'b1, 1'b0};
787: data_out = {8'd76, 8'd25, 1'b1, 1'b0};
788: data_out = {8'd77, 8'd25, 1'b1, 1'b0};
789: data_out = {8'd78, 8'd25, 1'b1, 1'b0};
790: data_out = {8'd85, 8'd25, 1'b1, 1'b0};
791: data_out = {8'd86, 8'd25, 1'b1, 1'b0};
792: data_out = {8'd87, 8'd25, 1'b1, 1'b0};
793: data_out = {8'd88, 8'd25, 1'b1, 1'b0};
794: data_out = {8'd89, 8'd25, 1'b1, 1'b0};
795: data_out = {8'd90, 8'd25, 1'b1, 1'b0};
796: data_out = {8'd97, 8'd25, 1'b1, 1'b0};
797: data_out = {8'd98, 8'd25, 1'b1, 1'b0};
798: data_out = {8'd99, 8'd25, 1'b1, 1'b0};
799: data_out = {8'd100, 8'd25, 1'b1, 1'b0};
800: data_out = {8'd101, 8'd25, 1'b1, 1'b0};
801: data_out = {8'd102, 8'd25, 1'b1, 1'b0};
802: data_out = {8'd116, 8'd25, 1'b1, 1'b0};
803: data_out = {8'd117, 8'd25, 1'b1, 1'b0};
804: data_out = {8'd118, 8'd25, 1'b1, 1'b0};
805: data_out = {8'd119, 8'd25, 1'b1, 1'b0};
806: data_out = {8'd120, 8'd25, 1'b1, 1'b0};
807: data_out = {8'd121, 8'd25, 1'b1, 1'b0};
808: data_out = {8'd127, 8'd25, 1'b1, 1'b0};
809: data_out = {8'd128, 8'd25, 1'b1, 1'b0};
810: data_out = {8'd129, 8'd25, 1'b1, 1'b0};
811: data_out = {8'd130, 8'd25, 1'b1, 1'b0};
812: data_out = {8'd131, 8'd25, 1'b1, 1'b0};
813: data_out = {8'd132, 8'd25, 1'b1, 1'b0};
814: data_out = {8'd146, 8'd25, 1'b1, 1'b0};
815: data_out = {8'd147, 8'd25, 1'b1, 1'b0};
816: data_out = {8'd148, 8'd25, 1'b1, 1'b0};
817: data_out = {8'd149, 8'd25, 1'b1, 1'b0};
818: data_out = {8'd150, 8'd25, 1'b1, 1'b0};
819: data_out = {8'd151, 8'd25, 1'b1, 1'b0};
820: data_out = {8'd187, 8'd25, 1'b1, 1'b0};
821: data_out = {8'd188, 8'd25, 1'b1, 1'b0};
822: data_out = {8'd189, 8'd25, 1'b1, 1'b0};
823: data_out = {8'd190, 8'd25, 1'b1, 1'b0};
824: data_out = {8'd191, 8'd25, 1'b1, 1'b0};
825: data_out = {8'd192, 8'd25, 1'b1, 1'b0};
826: data_out = {8'd206, 8'd25, 1'b1, 1'b0};
827: data_out = {8'd207, 8'd25, 1'b1, 1'b0};
828: data_out = {8'd208, 8'd25, 1'b1, 1'b0};
829: data_out = {8'd209, 8'd25, 1'b1, 1'b0};
830: data_out = {8'd210, 8'd25, 1'b1, 1'b0};
831: data_out = {8'd211, 8'd25, 1'b1, 1'b0};
832: data_out = {8'd6, 8'd26, 1'b1, 1'b0};
833: data_out = {8'd7, 8'd26, 1'b1, 1'b0};
834: data_out = {8'd8, 8'd26, 1'b1, 1'b0};
835: data_out = {8'd9, 8'd26, 1'b1, 1'b0};
836: data_out = {8'd10, 8'd26, 1'b1, 1'b0};
837: data_out = {8'd11, 8'd26, 1'b1, 1'b0};
838: data_out = {8'd25, 8'd26, 1'b1, 1'b0};
839: data_out = {8'd26, 8'd26, 1'b1, 1'b0};
840: data_out = {8'd27, 8'd26, 1'b1, 1'b0};
841: data_out = {8'd28, 8'd26, 1'b1, 1'b0};
842: data_out = {8'd29, 8'd26, 1'b1, 1'b0};
843: data_out = {8'd30, 8'd26, 1'b1, 1'b0};
844: data_out = {8'd36, 8'd26, 1'b1, 1'b0};
845: data_out = {8'd37, 8'd26, 1'b1, 1'b0};
846: data_out = {8'd38, 8'd26, 1'b1, 1'b0};
847: data_out = {8'd39, 8'd26, 1'b1, 1'b0};
848: data_out = {8'd40, 8'd26, 1'b1, 1'b0};
849: data_out = {8'd41, 8'd26, 1'b1, 1'b0};
850: data_out = {8'd55, 8'd26, 1'b1, 1'b0};
851: data_out = {8'd56, 8'd26, 1'b1, 1'b0};
852: data_out = {8'd57, 8'd26, 1'b1, 1'b0};
853: data_out = {8'd58, 8'd26, 1'b1, 1'b0};
854: data_out = {8'd59, 8'd26, 1'b1, 1'b0};
855: data_out = {8'd60, 8'd26, 1'b1, 1'b0};
856: data_out = {8'd73, 8'd26, 1'b1, 1'b0};
857: data_out = {8'd74, 8'd26, 1'b1, 1'b0};
858: data_out = {8'd75, 8'd26, 1'b1, 1'b0};
859: data_out = {8'd76, 8'd26, 1'b1, 1'b0};
860: data_out = {8'd77, 8'd26, 1'b1, 1'b0};
861: data_out = {8'd78, 8'd26, 1'b1, 1'b0};
862: data_out = {8'd85, 8'd26, 1'b1, 1'b0};
863: data_out = {8'd86, 8'd26, 1'b1, 1'b0};
864: data_out = {8'd87, 8'd26, 1'b1, 1'b0};
865: data_out = {8'd88, 8'd26, 1'b1, 1'b0};
866: data_out = {8'd89, 8'd26, 1'b1, 1'b0};
867: data_out = {8'd90, 8'd26, 1'b1, 1'b0};
868: data_out = {8'd97, 8'd26, 1'b1, 1'b0};
869: data_out = {8'd98, 8'd26, 1'b1, 1'b0};
870: data_out = {8'd99, 8'd26, 1'b1, 1'b0};
871: data_out = {8'd100, 8'd26, 1'b1, 1'b0};
872: data_out = {8'd101, 8'd26, 1'b1, 1'b0};
873: data_out = {8'd102, 8'd26, 1'b1, 1'b0};
874: data_out = {8'd116, 8'd26, 1'b1, 1'b0};
875: data_out = {8'd117, 8'd26, 1'b1, 1'b0};
876: data_out = {8'd118, 8'd26, 1'b1, 1'b0};
877: data_out = {8'd119, 8'd26, 1'b1, 1'b0};
878: data_out = {8'd120, 8'd26, 1'b1, 1'b0};
879: data_out = {8'd121, 8'd26, 1'b1, 1'b0};
880: data_out = {8'd127, 8'd26, 1'b1, 1'b0};
881: data_out = {8'd128, 8'd26, 1'b1, 1'b0};
882: data_out = {8'd129, 8'd26, 1'b1, 1'b0};
883: data_out = {8'd130, 8'd26, 1'b1, 1'b0};
884: data_out = {8'd131, 8'd26, 1'b1, 1'b0};
885: data_out = {8'd132, 8'd26, 1'b1, 1'b0};
886: data_out = {8'd146, 8'd26, 1'b1, 1'b0};
887: data_out = {8'd147, 8'd26, 1'b1, 1'b0};
888: data_out = {8'd148, 8'd26, 1'b1, 1'b0};
889: data_out = {8'd149, 8'd26, 1'b1, 1'b0};
890: data_out = {8'd150, 8'd26, 1'b1, 1'b0};
891: data_out = {8'd151, 8'd26, 1'b1, 1'b0};
892: data_out = {8'd187, 8'd26, 1'b1, 1'b0};
893: data_out = {8'd188, 8'd26, 1'b1, 1'b0};
894: data_out = {8'd189, 8'd26, 1'b1, 1'b0};
895: data_out = {8'd190, 8'd26, 1'b1, 1'b0};
896: data_out = {8'd191, 8'd26, 1'b1, 1'b0};
897: data_out = {8'd192, 8'd26, 1'b1, 1'b0};
898: data_out = {8'd206, 8'd26, 1'b1, 1'b0};
899: data_out = {8'd207, 8'd26, 1'b1, 1'b0};
900: data_out = {8'd208, 8'd26, 1'b1, 1'b0};
901: data_out = {8'd209, 8'd26, 1'b1, 1'b0};
902: data_out = {8'd210, 8'd26, 1'b1, 1'b0};
903: data_out = {8'd211, 8'd26, 1'b1, 1'b0};
904: data_out = {8'd6, 8'd27, 1'b1, 1'b0};
905: data_out = {8'd7, 8'd27, 1'b1, 1'b0};
906: data_out = {8'd8, 8'd27, 1'b1, 1'b0};
907: data_out = {8'd9, 8'd27, 1'b1, 1'b0};
908: data_out = {8'd10, 8'd27, 1'b1, 1'b0};
909: data_out = {8'd11, 8'd27, 1'b1, 1'b0};
910: data_out = {8'd25, 8'd27, 1'b1, 1'b0};
911: data_out = {8'd26, 8'd27, 1'b1, 1'b0};
912: data_out = {8'd27, 8'd27, 1'b1, 1'b0};
913: data_out = {8'd28, 8'd27, 1'b1, 1'b0};
914: data_out = {8'd29, 8'd27, 1'b1, 1'b0};
915: data_out = {8'd30, 8'd27, 1'b1, 1'b0};
916: data_out = {8'd36, 8'd27, 1'b1, 1'b0};
917: data_out = {8'd37, 8'd27, 1'b1, 1'b0};
918: data_out = {8'd38, 8'd27, 1'b1, 1'b0};
919: data_out = {8'd39, 8'd27, 1'b1, 1'b0};
920: data_out = {8'd40, 8'd27, 1'b1, 1'b0};
921: data_out = {8'd41, 8'd27, 1'b1, 1'b0};
922: data_out = {8'd55, 8'd27, 1'b1, 1'b0};
923: data_out = {8'd56, 8'd27, 1'b1, 1'b0};
924: data_out = {8'd57, 8'd27, 1'b1, 1'b0};
925: data_out = {8'd58, 8'd27, 1'b1, 1'b0};
926: data_out = {8'd59, 8'd27, 1'b1, 1'b0};
927: data_out = {8'd60, 8'd27, 1'b1, 1'b0};
928: data_out = {8'd73, 8'd27, 1'b1, 1'b0};
929: data_out = {8'd74, 8'd27, 1'b1, 1'b0};
930: data_out = {8'd75, 8'd27, 1'b1, 1'b0};
931: data_out = {8'd76, 8'd27, 1'b1, 1'b0};
932: data_out = {8'd77, 8'd27, 1'b1, 1'b0};
933: data_out = {8'd78, 8'd27, 1'b1, 1'b0};
934: data_out = {8'd85, 8'd27, 1'b1, 1'b0};
935: data_out = {8'd86, 8'd27, 1'b1, 1'b0};
936: data_out = {8'd87, 8'd27, 1'b1, 1'b0};
937: data_out = {8'd88, 8'd27, 1'b1, 1'b0};
938: data_out = {8'd89, 8'd27, 1'b1, 1'b0};
939: data_out = {8'd90, 8'd27, 1'b1, 1'b0};
940: data_out = {8'd97, 8'd27, 1'b1, 1'b0};
941: data_out = {8'd98, 8'd27, 1'b1, 1'b0};
942: data_out = {8'd99, 8'd27, 1'b1, 1'b0};
943: data_out = {8'd100, 8'd27, 1'b1, 1'b0};
944: data_out = {8'd101, 8'd27, 1'b1, 1'b0};
945: data_out = {8'd102, 8'd27, 1'b1, 1'b0};
946: data_out = {8'd116, 8'd27, 1'b1, 1'b0};
947: data_out = {8'd117, 8'd27, 1'b1, 1'b0};
948: data_out = {8'd118, 8'd27, 1'b1, 1'b0};
949: data_out = {8'd119, 8'd27, 1'b1, 1'b0};
950: data_out = {8'd120, 8'd27, 1'b1, 1'b0};
951: data_out = {8'd121, 8'd27, 1'b1, 1'b0};
952: data_out = {8'd127, 8'd27, 1'b1, 1'b0};
953: data_out = {8'd128, 8'd27, 1'b1, 1'b0};
954: data_out = {8'd129, 8'd27, 1'b1, 1'b0};
955: data_out = {8'd130, 8'd27, 1'b1, 1'b0};
956: data_out = {8'd131, 8'd27, 1'b1, 1'b0};
957: data_out = {8'd132, 8'd27, 1'b1, 1'b0};
958: data_out = {8'd146, 8'd27, 1'b1, 1'b0};
959: data_out = {8'd147, 8'd27, 1'b1, 1'b0};
960: data_out = {8'd148, 8'd27, 1'b1, 1'b0};
961: data_out = {8'd149, 8'd27, 1'b1, 1'b0};
962: data_out = {8'd150, 8'd27, 1'b1, 1'b0};
963: data_out = {8'd151, 8'd27, 1'b1, 1'b0};
964: data_out = {8'd187, 8'd27, 1'b1, 1'b0};
965: data_out = {8'd188, 8'd27, 1'b1, 1'b0};
966: data_out = {8'd189, 8'd27, 1'b1, 1'b0};
967: data_out = {8'd190, 8'd27, 1'b1, 1'b0};
968: data_out = {8'd191, 8'd27, 1'b1, 1'b0};
969: data_out = {8'd192, 8'd27, 1'b1, 1'b0};
970: data_out = {8'd206, 8'd27, 1'b1, 1'b0};
971: data_out = {8'd207, 8'd27, 1'b1, 1'b0};
972: data_out = {8'd208, 8'd27, 1'b1, 1'b0};
973: data_out = {8'd209, 8'd27, 1'b1, 1'b0};
974: data_out = {8'd210, 8'd27, 1'b1, 1'b0};
975: data_out = {8'd211, 8'd27, 1'b1, 1'b0};
976: data_out = {8'd6, 8'd28, 1'b1, 1'b0};
977: data_out = {8'd7, 8'd28, 1'b1, 1'b0};
978: data_out = {8'd8, 8'd28, 1'b1, 1'b0};
979: data_out = {8'd9, 8'd28, 1'b1, 1'b0};
980: data_out = {8'd10, 8'd28, 1'b1, 1'b0};
981: data_out = {8'd11, 8'd28, 1'b1, 1'b0};
982: data_out = {8'd25, 8'd28, 1'b1, 1'b0};
983: data_out = {8'd26, 8'd28, 1'b1, 1'b0};
984: data_out = {8'd27, 8'd28, 1'b1, 1'b0};
985: data_out = {8'd28, 8'd28, 1'b1, 1'b0};
986: data_out = {8'd29, 8'd28, 1'b1, 1'b0};
987: data_out = {8'd30, 8'd28, 1'b1, 1'b0};
988: data_out = {8'd36, 8'd28, 1'b1, 1'b0};
989: data_out = {8'd37, 8'd28, 1'b1, 1'b0};
990: data_out = {8'd38, 8'd28, 1'b1, 1'b0};
991: data_out = {8'd39, 8'd28, 1'b1, 1'b0};
992: data_out = {8'd40, 8'd28, 1'b1, 1'b0};
993: data_out = {8'd41, 8'd28, 1'b1, 1'b0};
994: data_out = {8'd55, 8'd28, 1'b1, 1'b0};
995: data_out = {8'd56, 8'd28, 1'b1, 1'b0};
996: data_out = {8'd57, 8'd28, 1'b1, 1'b0};
997: data_out = {8'd58, 8'd28, 1'b1, 1'b0};
998: data_out = {8'd59, 8'd28, 1'b1, 1'b0};
999: data_out = {8'd60, 8'd28, 1'b1, 1'b0};
1000: data_out = {8'd73, 8'd28, 1'b1, 1'b0};
1001: data_out = {8'd74, 8'd28, 1'b1, 1'b0};
1002: data_out = {8'd75, 8'd28, 1'b1, 1'b0};
1003: data_out = {8'd76, 8'd28, 1'b1, 1'b0};
1004: data_out = {8'd77, 8'd28, 1'b1, 1'b0};
1005: data_out = {8'd78, 8'd28, 1'b1, 1'b0};
1006: data_out = {8'd85, 8'd28, 1'b1, 1'b0};
1007: data_out = {8'd86, 8'd28, 1'b1, 1'b0};
1008: data_out = {8'd87, 8'd28, 1'b1, 1'b0};
1009: data_out = {8'd88, 8'd28, 1'b1, 1'b0};
1010: data_out = {8'd89, 8'd28, 1'b1, 1'b0};
1011: data_out = {8'd90, 8'd28, 1'b1, 1'b0};
1012: data_out = {8'd97, 8'd28, 1'b1, 1'b0};
1013: data_out = {8'd98, 8'd28, 1'b1, 1'b0};
1014: data_out = {8'd99, 8'd28, 1'b1, 1'b0};
1015: data_out = {8'd100, 8'd28, 1'b1, 1'b0};
1016: data_out = {8'd101, 8'd28, 1'b1, 1'b0};
1017: data_out = {8'd102, 8'd28, 1'b1, 1'b0};
1018: data_out = {8'd116, 8'd28, 1'b1, 1'b0};
1019: data_out = {8'd117, 8'd28, 1'b1, 1'b0};
1020: data_out = {8'd118, 8'd28, 1'b1, 1'b0};
1021: data_out = {8'd119, 8'd28, 1'b1, 1'b0};
1022: data_out = {8'd120, 8'd28, 1'b1, 1'b0};
1023: data_out = {8'd121, 8'd28, 1'b1, 1'b0};
1024: data_out = {8'd127, 8'd28, 1'b1, 1'b0};
1025: data_out = {8'd128, 8'd28, 1'b1, 1'b0};
1026: data_out = {8'd129, 8'd28, 1'b1, 1'b0};
1027: data_out = {8'd130, 8'd28, 1'b1, 1'b0};
1028: data_out = {8'd131, 8'd28, 1'b1, 1'b0};
1029: data_out = {8'd132, 8'd28, 1'b1, 1'b0};
1030: data_out = {8'd146, 8'd28, 1'b1, 1'b0};
1031: data_out = {8'd147, 8'd28, 1'b1, 1'b0};
1032: data_out = {8'd148, 8'd28, 1'b1, 1'b0};
1033: data_out = {8'd149, 8'd28, 1'b1, 1'b0};
1034: data_out = {8'd150, 8'd28, 1'b1, 1'b0};
1035: data_out = {8'd151, 8'd28, 1'b1, 1'b0};
1036: data_out = {8'd187, 8'd28, 1'b1, 1'b0};
1037: data_out = {8'd188, 8'd28, 1'b1, 1'b0};
1038: data_out = {8'd189, 8'd28, 1'b1, 1'b0};
1039: data_out = {8'd190, 8'd28, 1'b1, 1'b0};
1040: data_out = {8'd191, 8'd28, 1'b1, 1'b0};
1041: data_out = {8'd192, 8'd28, 1'b1, 1'b0};
1042: data_out = {8'd206, 8'd28, 1'b1, 1'b0};
1043: data_out = {8'd207, 8'd28, 1'b1, 1'b0};
1044: data_out = {8'd208, 8'd28, 1'b1, 1'b0};
1045: data_out = {8'd209, 8'd28, 1'b1, 1'b0};
1046: data_out = {8'd210, 8'd28, 1'b1, 1'b0};
1047: data_out = {8'd211, 8'd28, 1'b1, 1'b0};
1048: data_out = {8'd6, 8'd29, 1'b1, 1'b0};
1049: data_out = {8'd7, 8'd29, 1'b1, 1'b0};
1050: data_out = {8'd8, 8'd29, 1'b1, 1'b0};
1051: data_out = {8'd9, 8'd29, 1'b1, 1'b0};
1052: data_out = {8'd10, 8'd29, 1'b1, 1'b0};
1053: data_out = {8'd11, 8'd29, 1'b1, 1'b0};
1054: data_out = {8'd25, 8'd29, 1'b1, 1'b0};
1055: data_out = {8'd26, 8'd29, 1'b1, 1'b0};
1056: data_out = {8'd27, 8'd29, 1'b1, 1'b0};
1057: data_out = {8'd28, 8'd29, 1'b1, 1'b0};
1058: data_out = {8'd29, 8'd29, 1'b1, 1'b0};
1059: data_out = {8'd30, 8'd29, 1'b1, 1'b0};
1060: data_out = {8'd36, 8'd29, 1'b1, 1'b0};
1061: data_out = {8'd37, 8'd29, 1'b1, 1'b0};
1062: data_out = {8'd38, 8'd29, 1'b1, 1'b0};
1063: data_out = {8'd39, 8'd29, 1'b1, 1'b0};
1064: data_out = {8'd40, 8'd29, 1'b1, 1'b0};
1065: data_out = {8'd41, 8'd29, 1'b1, 1'b0};
1066: data_out = {8'd55, 8'd29, 1'b1, 1'b0};
1067: data_out = {8'd56, 8'd29, 1'b1, 1'b0};
1068: data_out = {8'd57, 8'd29, 1'b1, 1'b0};
1069: data_out = {8'd58, 8'd29, 1'b1, 1'b0};
1070: data_out = {8'd59, 8'd29, 1'b1, 1'b0};
1071: data_out = {8'd60, 8'd29, 1'b1, 1'b0};
1072: data_out = {8'd73, 8'd29, 1'b1, 1'b0};
1073: data_out = {8'd74, 8'd29, 1'b1, 1'b0};
1074: data_out = {8'd75, 8'd29, 1'b1, 1'b0};
1075: data_out = {8'd76, 8'd29, 1'b1, 1'b0};
1076: data_out = {8'd77, 8'd29, 1'b1, 1'b0};
1077: data_out = {8'd78, 8'd29, 1'b1, 1'b0};
1078: data_out = {8'd85, 8'd29, 1'b1, 1'b0};
1079: data_out = {8'd86, 8'd29, 1'b1, 1'b0};
1080: data_out = {8'd87, 8'd29, 1'b1, 1'b0};
1081: data_out = {8'd88, 8'd29, 1'b1, 1'b0};
1082: data_out = {8'd89, 8'd29, 1'b1, 1'b0};
1083: data_out = {8'd90, 8'd29, 1'b1, 1'b0};
1084: data_out = {8'd97, 8'd29, 1'b1, 1'b0};
1085: data_out = {8'd98, 8'd29, 1'b1, 1'b0};
1086: data_out = {8'd99, 8'd29, 1'b1, 1'b0};
1087: data_out = {8'd100, 8'd29, 1'b1, 1'b0};
1088: data_out = {8'd101, 8'd29, 1'b1, 1'b0};
1089: data_out = {8'd102, 8'd29, 1'b1, 1'b0};
1090: data_out = {8'd116, 8'd29, 1'b1, 1'b0};
1091: data_out = {8'd117, 8'd29, 1'b1, 1'b0};
1092: data_out = {8'd118, 8'd29, 1'b1, 1'b0};
1093: data_out = {8'd119, 8'd29, 1'b1, 1'b0};
1094: data_out = {8'd120, 8'd29, 1'b1, 1'b0};
1095: data_out = {8'd121, 8'd29, 1'b1, 1'b0};
1096: data_out = {8'd127, 8'd29, 1'b1, 1'b0};
1097: data_out = {8'd128, 8'd29, 1'b1, 1'b0};
1098: data_out = {8'd129, 8'd29, 1'b1, 1'b0};
1099: data_out = {8'd130, 8'd29, 1'b1, 1'b0};
1100: data_out = {8'd131, 8'd29, 1'b1, 1'b0};
1101: data_out = {8'd132, 8'd29, 1'b1, 1'b0};
1102: data_out = {8'd146, 8'd29, 1'b1, 1'b0};
1103: data_out = {8'd147, 8'd29, 1'b1, 1'b0};
1104: data_out = {8'd148, 8'd29, 1'b1, 1'b0};
1105: data_out = {8'd149, 8'd29, 1'b1, 1'b0};
1106: data_out = {8'd150, 8'd29, 1'b1, 1'b0};
1107: data_out = {8'd151, 8'd29, 1'b1, 1'b0};
1108: data_out = {8'd187, 8'd29, 1'b1, 1'b0};
1109: data_out = {8'd188, 8'd29, 1'b1, 1'b0};
1110: data_out = {8'd189, 8'd29, 1'b1, 1'b0};
1111: data_out = {8'd190, 8'd29, 1'b1, 1'b0};
1112: data_out = {8'd191, 8'd29, 1'b1, 1'b0};
1113: data_out = {8'd192, 8'd29, 1'b1, 1'b0};
1114: data_out = {8'd206, 8'd29, 1'b1, 1'b0};
1115: data_out = {8'd207, 8'd29, 1'b1, 1'b0};
1116: data_out = {8'd208, 8'd29, 1'b1, 1'b0};
1117: data_out = {8'd209, 8'd29, 1'b1, 1'b0};
1118: data_out = {8'd210, 8'd29, 1'b1, 1'b0};
1119: data_out = {8'd211, 8'd29, 1'b1, 1'b0};
1120: data_out = {8'd6, 8'd30, 1'b1, 1'b0};
1121: data_out = {8'd7, 8'd30, 1'b1, 1'b0};
1122: data_out = {8'd8, 8'd30, 1'b1, 1'b0};
1123: data_out = {8'd9, 8'd30, 1'b1, 1'b0};
1124: data_out = {8'd10, 8'd30, 1'b1, 1'b0};
1125: data_out = {8'd11, 8'd30, 1'b1, 1'b0};
1126: data_out = {8'd25, 8'd30, 1'b1, 1'b0};
1127: data_out = {8'd26, 8'd30, 1'b1, 1'b0};
1128: data_out = {8'd27, 8'd30, 1'b1, 1'b0};
1129: data_out = {8'd28, 8'd30, 1'b1, 1'b0};
1130: data_out = {8'd29, 8'd30, 1'b1, 1'b0};
1131: data_out = {8'd30, 8'd30, 1'b1, 1'b0};
1132: data_out = {8'd36, 8'd30, 1'b1, 1'b0};
1133: data_out = {8'd37, 8'd30, 1'b1, 1'b0};
1134: data_out = {8'd38, 8'd30, 1'b1, 1'b0};
1135: data_out = {8'd39, 8'd30, 1'b1, 1'b0};
1136: data_out = {8'd40, 8'd30, 1'b1, 1'b0};
1137: data_out = {8'd41, 8'd30, 1'b1, 1'b0};
1138: data_out = {8'd55, 8'd30, 1'b1, 1'b0};
1139: data_out = {8'd56, 8'd30, 1'b1, 1'b0};
1140: data_out = {8'd57, 8'd30, 1'b1, 1'b0};
1141: data_out = {8'd58, 8'd30, 1'b1, 1'b0};
1142: data_out = {8'd59, 8'd30, 1'b1, 1'b0};
1143: data_out = {8'd60, 8'd30, 1'b1, 1'b0};
1144: data_out = {8'd73, 8'd30, 1'b1, 1'b0};
1145: data_out = {8'd74, 8'd30, 1'b1, 1'b0};
1146: data_out = {8'd75, 8'd30, 1'b1, 1'b0};
1147: data_out = {8'd76, 8'd30, 1'b1, 1'b0};
1148: data_out = {8'd77, 8'd30, 1'b1, 1'b0};
1149: data_out = {8'd78, 8'd30, 1'b1, 1'b0};
1150: data_out = {8'd85, 8'd30, 1'b1, 1'b0};
1151: data_out = {8'd86, 8'd30, 1'b1, 1'b0};
1152: data_out = {8'd87, 8'd30, 1'b1, 1'b0};
1153: data_out = {8'd88, 8'd30, 1'b1, 1'b0};
1154: data_out = {8'd89, 8'd30, 1'b1, 1'b0};
1155: data_out = {8'd90, 8'd30, 1'b1, 1'b0};
1156: data_out = {8'd97, 8'd30, 1'b1, 1'b0};
1157: data_out = {8'd98, 8'd30, 1'b1, 1'b0};
1158: data_out = {8'd99, 8'd30, 1'b1, 1'b0};
1159: data_out = {8'd100, 8'd30, 1'b1, 1'b0};
1160: data_out = {8'd101, 8'd30, 1'b1, 1'b0};
1161: data_out = {8'd102, 8'd30, 1'b1, 1'b0};
1162: data_out = {8'd116, 8'd30, 1'b1, 1'b0};
1163: data_out = {8'd117, 8'd30, 1'b1, 1'b0};
1164: data_out = {8'd118, 8'd30, 1'b1, 1'b0};
1165: data_out = {8'd119, 8'd30, 1'b1, 1'b0};
1166: data_out = {8'd120, 8'd30, 1'b1, 1'b0};
1167: data_out = {8'd121, 8'd30, 1'b1, 1'b0};
1168: data_out = {8'd127, 8'd30, 1'b1, 1'b0};
1169: data_out = {8'd128, 8'd30, 1'b1, 1'b0};
1170: data_out = {8'd129, 8'd30, 1'b1, 1'b0};
1171: data_out = {8'd130, 8'd30, 1'b1, 1'b0};
1172: data_out = {8'd131, 8'd30, 1'b1, 1'b0};
1173: data_out = {8'd132, 8'd30, 1'b1, 1'b0};
1174: data_out = {8'd146, 8'd30, 1'b1, 1'b0};
1175: data_out = {8'd147, 8'd30, 1'b1, 1'b0};
1176: data_out = {8'd148, 8'd30, 1'b1, 1'b0};
1177: data_out = {8'd149, 8'd30, 1'b1, 1'b0};
1178: data_out = {8'd150, 8'd30, 1'b1, 1'b0};
1179: data_out = {8'd151, 8'd30, 1'b1, 1'b0};
1180: data_out = {8'd187, 8'd30, 1'b1, 1'b0};
1181: data_out = {8'd188, 8'd30, 1'b1, 1'b0};
1182: data_out = {8'd189, 8'd30, 1'b1, 1'b0};
1183: data_out = {8'd190, 8'd30, 1'b1, 1'b0};
1184: data_out = {8'd191, 8'd30, 1'b1, 1'b0};
1185: data_out = {8'd192, 8'd30, 1'b1, 1'b0};
1186: data_out = {8'd206, 8'd30, 1'b1, 1'b0};
1187: data_out = {8'd207, 8'd30, 1'b1, 1'b0};
1188: data_out = {8'd208, 8'd30, 1'b1, 1'b0};
1189: data_out = {8'd209, 8'd30, 1'b1, 1'b0};
1190: data_out = {8'd210, 8'd30, 1'b1, 1'b0};
1191: data_out = {8'd211, 8'd30, 1'b1, 1'b0};
1192: data_out = {8'd6, 8'd31, 1'b1, 1'b0};
1193: data_out = {8'd7, 8'd31, 1'b1, 1'b0};
1194: data_out = {8'd8, 8'd31, 1'b1, 1'b0};
1195: data_out = {8'd9, 8'd31, 1'b1, 1'b0};
1196: data_out = {8'd10, 8'd31, 1'b1, 1'b0};
1197: data_out = {8'd11, 8'd31, 1'b1, 1'b0};
1198: data_out = {8'd25, 8'd31, 1'b1, 1'b0};
1199: data_out = {8'd26, 8'd31, 1'b1, 1'b0};
1200: data_out = {8'd27, 8'd31, 1'b1, 1'b0};
1201: data_out = {8'd28, 8'd31, 1'b1, 1'b0};
1202: data_out = {8'd29, 8'd31, 1'b1, 1'b0};
1203: data_out = {8'd30, 8'd31, 1'b1, 1'b0};
1204: data_out = {8'd36, 8'd31, 1'b1, 1'b0};
1205: data_out = {8'd37, 8'd31, 1'b1, 1'b0};
1206: data_out = {8'd38, 8'd31, 1'b1, 1'b0};
1207: data_out = {8'd39, 8'd31, 1'b1, 1'b0};
1208: data_out = {8'd40, 8'd31, 1'b1, 1'b0};
1209: data_out = {8'd41, 8'd31, 1'b1, 1'b0};
1210: data_out = {8'd55, 8'd31, 1'b1, 1'b0};
1211: data_out = {8'd56, 8'd31, 1'b1, 1'b0};
1212: data_out = {8'd57, 8'd31, 1'b1, 1'b0};
1213: data_out = {8'd58, 8'd31, 1'b1, 1'b0};
1214: data_out = {8'd59, 8'd31, 1'b1, 1'b0};
1215: data_out = {8'd60, 8'd31, 1'b1, 1'b0};
1216: data_out = {8'd73, 8'd31, 1'b1, 1'b0};
1217: data_out = {8'd74, 8'd31, 1'b1, 1'b0};
1218: data_out = {8'd75, 8'd31, 1'b1, 1'b0};
1219: data_out = {8'd76, 8'd31, 1'b1, 1'b0};
1220: data_out = {8'd77, 8'd31, 1'b1, 1'b0};
1221: data_out = {8'd78, 8'd31, 1'b1, 1'b0};
1222: data_out = {8'd116, 8'd31, 1'b1, 1'b0};
1223: data_out = {8'd117, 8'd31, 1'b1, 1'b0};
1224: data_out = {8'd118, 8'd31, 1'b1, 1'b0};
1225: data_out = {8'd119, 8'd31, 1'b1, 1'b0};
1226: data_out = {8'd120, 8'd31, 1'b1, 1'b0};
1227: data_out = {8'd121, 8'd31, 1'b1, 1'b0};
1228: data_out = {8'd127, 8'd31, 1'b1, 1'b0};
1229: data_out = {8'd128, 8'd31, 1'b1, 1'b0};
1230: data_out = {8'd129, 8'd31, 1'b1, 1'b0};
1231: data_out = {8'd130, 8'd31, 1'b1, 1'b0};
1232: data_out = {8'd131, 8'd31, 1'b1, 1'b0};
1233: data_out = {8'd132, 8'd31, 1'b1, 1'b0};
1234: data_out = {8'd146, 8'd31, 1'b1, 1'b0};
1235: data_out = {8'd147, 8'd31, 1'b1, 1'b0};
1236: data_out = {8'd148, 8'd31, 1'b1, 1'b0};
1237: data_out = {8'd149, 8'd31, 1'b1, 1'b0};
1238: data_out = {8'd150, 8'd31, 1'b1, 1'b0};
1239: data_out = {8'd151, 8'd31, 1'b1, 1'b0};
1240: data_out = {8'd206, 8'd31, 1'b1, 1'b0};
1241: data_out = {8'd207, 8'd31, 1'b1, 1'b0};
1242: data_out = {8'd208, 8'd31, 1'b1, 1'b0};
1243: data_out = {8'd209, 8'd31, 1'b1, 1'b0};
1244: data_out = {8'd210, 8'd31, 1'b1, 1'b0};
1245: data_out = {8'd211, 8'd31, 1'b1, 1'b0};
1246: data_out = {8'd6, 8'd32, 1'b1, 1'b0};
1247: data_out = {8'd7, 8'd32, 1'b1, 1'b0};
1248: data_out = {8'd8, 8'd32, 1'b1, 1'b0};
1249: data_out = {8'd9, 8'd32, 1'b1, 1'b0};
1250: data_out = {8'd10, 8'd32, 1'b1, 1'b0};
1251: data_out = {8'd11, 8'd32, 1'b1, 1'b0};
1252: data_out = {8'd25, 8'd32, 1'b1, 1'b0};
1253: data_out = {8'd26, 8'd32, 1'b1, 1'b0};
1254: data_out = {8'd27, 8'd32, 1'b1, 1'b0};
1255: data_out = {8'd28, 8'd32, 1'b1, 1'b0};
1256: data_out = {8'd29, 8'd32, 1'b1, 1'b0};
1257: data_out = {8'd30, 8'd32, 1'b1, 1'b0};
1258: data_out = {8'd36, 8'd32, 1'b1, 1'b0};
1259: data_out = {8'd37, 8'd32, 1'b1, 1'b0};
1260: data_out = {8'd38, 8'd32, 1'b1, 1'b0};
1261: data_out = {8'd39, 8'd32, 1'b1, 1'b0};
1262: data_out = {8'd40, 8'd32, 1'b1, 1'b0};
1263: data_out = {8'd41, 8'd32, 1'b1, 1'b0};
1264: data_out = {8'd55, 8'd32, 1'b1, 1'b0};
1265: data_out = {8'd56, 8'd32, 1'b1, 1'b0};
1266: data_out = {8'd57, 8'd32, 1'b1, 1'b0};
1267: data_out = {8'd58, 8'd32, 1'b1, 1'b0};
1268: data_out = {8'd59, 8'd32, 1'b1, 1'b0};
1269: data_out = {8'd60, 8'd32, 1'b1, 1'b0};
1270: data_out = {8'd73, 8'd32, 1'b1, 1'b0};
1271: data_out = {8'd74, 8'd32, 1'b1, 1'b0};
1272: data_out = {8'd75, 8'd32, 1'b1, 1'b0};
1273: data_out = {8'd76, 8'd32, 1'b1, 1'b0};
1274: data_out = {8'd77, 8'd32, 1'b1, 1'b0};
1275: data_out = {8'd78, 8'd32, 1'b1, 1'b0};
1276: data_out = {8'd116, 8'd32, 1'b1, 1'b0};
1277: data_out = {8'd117, 8'd32, 1'b1, 1'b0};
1278: data_out = {8'd118, 8'd32, 1'b1, 1'b0};
1279: data_out = {8'd119, 8'd32, 1'b1, 1'b0};
1280: data_out = {8'd120, 8'd32, 1'b1, 1'b0};
1281: data_out = {8'd121, 8'd32, 1'b1, 1'b0};
1282: data_out = {8'd127, 8'd32, 1'b1, 1'b0};
1283: data_out = {8'd128, 8'd32, 1'b1, 1'b0};
1284: data_out = {8'd129, 8'd32, 1'b1, 1'b0};
1285: data_out = {8'd130, 8'd32, 1'b1, 1'b0};
1286: data_out = {8'd131, 8'd32, 1'b1, 1'b0};
1287: data_out = {8'd132, 8'd32, 1'b1, 1'b0};
1288: data_out = {8'd146, 8'd32, 1'b1, 1'b0};
1289: data_out = {8'd147, 8'd32, 1'b1, 1'b0};
1290: data_out = {8'd148, 8'd32, 1'b1, 1'b0};
1291: data_out = {8'd149, 8'd32, 1'b1, 1'b0};
1292: data_out = {8'd150, 8'd32, 1'b1, 1'b0};
1293: data_out = {8'd151, 8'd32, 1'b1, 1'b0};
1294: data_out = {8'd206, 8'd32, 1'b1, 1'b0};
1295: data_out = {8'd207, 8'd32, 1'b1, 1'b0};
1296: data_out = {8'd208, 8'd32, 1'b1, 1'b0};
1297: data_out = {8'd209, 8'd32, 1'b1, 1'b0};
1298: data_out = {8'd210, 8'd32, 1'b1, 1'b0};
1299: data_out = {8'd211, 8'd32, 1'b1, 1'b0};
1300: data_out = {8'd6, 8'd33, 1'b1, 1'b0};
1301: data_out = {8'd7, 8'd33, 1'b1, 1'b0};
1302: data_out = {8'd8, 8'd33, 1'b1, 1'b0};
1303: data_out = {8'd9, 8'd33, 1'b1, 1'b0};
1304: data_out = {8'd10, 8'd33, 1'b1, 1'b0};
1305: data_out = {8'd11, 8'd33, 1'b1, 1'b0};
1306: data_out = {8'd25, 8'd33, 1'b1, 1'b0};
1307: data_out = {8'd26, 8'd33, 1'b1, 1'b0};
1308: data_out = {8'd27, 8'd33, 1'b1, 1'b0};
1309: data_out = {8'd28, 8'd33, 1'b1, 1'b0};
1310: data_out = {8'd29, 8'd33, 1'b1, 1'b0};
1311: data_out = {8'd30, 8'd33, 1'b1, 1'b0};
1312: data_out = {8'd36, 8'd33, 1'b1, 1'b0};
1313: data_out = {8'd37, 8'd33, 1'b1, 1'b0};
1314: data_out = {8'd38, 8'd33, 1'b1, 1'b0};
1315: data_out = {8'd39, 8'd33, 1'b1, 1'b0};
1316: data_out = {8'd40, 8'd33, 1'b1, 1'b0};
1317: data_out = {8'd41, 8'd33, 1'b1, 1'b0};
1318: data_out = {8'd55, 8'd33, 1'b1, 1'b0};
1319: data_out = {8'd56, 8'd33, 1'b1, 1'b0};
1320: data_out = {8'd57, 8'd33, 1'b1, 1'b0};
1321: data_out = {8'd58, 8'd33, 1'b1, 1'b0};
1322: data_out = {8'd59, 8'd33, 1'b1, 1'b0};
1323: data_out = {8'd60, 8'd33, 1'b1, 1'b0};
1324: data_out = {8'd73, 8'd33, 1'b1, 1'b0};
1325: data_out = {8'd74, 8'd33, 1'b1, 1'b0};
1326: data_out = {8'd75, 8'd33, 1'b1, 1'b0};
1327: data_out = {8'd76, 8'd33, 1'b1, 1'b0};
1328: data_out = {8'd77, 8'd33, 1'b1, 1'b0};
1329: data_out = {8'd78, 8'd33, 1'b1, 1'b0};
1330: data_out = {8'd113, 8'd33, 1'b1, 1'b0};
1331: data_out = {8'd114, 8'd33, 1'b1, 1'b0};
1332: data_out = {8'd115, 8'd33, 1'b1, 1'b0};
1333: data_out = {8'd116, 8'd33, 1'b1, 1'b0};
1334: data_out = {8'd117, 8'd33, 1'b1, 1'b0};
1335: data_out = {8'd118, 8'd33, 1'b1, 1'b0};
1336: data_out = {8'd119, 8'd33, 1'b1, 1'b0};
1337: data_out = {8'd120, 8'd33, 1'b1, 1'b0};
1338: data_out = {8'd121, 8'd33, 1'b1, 1'b0};
1339: data_out = {8'd127, 8'd33, 1'b1, 1'b0};
1340: data_out = {8'd128, 8'd33, 1'b1, 1'b0};
1341: data_out = {8'd129, 8'd33, 1'b1, 1'b0};
1342: data_out = {8'd130, 8'd33, 1'b1, 1'b0};
1343: data_out = {8'd131, 8'd33, 1'b1, 1'b0};
1344: data_out = {8'd132, 8'd33, 1'b1, 1'b0};
1345: data_out = {8'd146, 8'd33, 1'b1, 1'b0};
1346: data_out = {8'd147, 8'd33, 1'b1, 1'b0};
1347: data_out = {8'd148, 8'd33, 1'b1, 1'b0};
1348: data_out = {8'd149, 8'd33, 1'b1, 1'b0};
1349: data_out = {8'd150, 8'd33, 1'b1, 1'b0};
1350: data_out = {8'd151, 8'd33, 1'b1, 1'b0};
1351: data_out = {8'd203, 8'd33, 1'b1, 1'b0};
1352: data_out = {8'd204, 8'd33, 1'b1, 1'b0};
1353: data_out = {8'd205, 8'd33, 1'b1, 1'b0};
1354: data_out = {8'd206, 8'd33, 1'b1, 1'b0};
1355: data_out = {8'd207, 8'd33, 1'b1, 1'b0};
1356: data_out = {8'd208, 8'd33, 1'b1, 1'b0};
1357: data_out = {8'd209, 8'd33, 1'b1, 1'b0};
1358: data_out = {8'd210, 8'd33, 1'b1, 1'b0};
1359: data_out = {8'd211, 8'd33, 1'b1, 1'b0};
1360: data_out = {8'd6, 8'd34, 1'b1, 1'b0};
1361: data_out = {8'd7, 8'd34, 1'b1, 1'b0};
1362: data_out = {8'd8, 8'd34, 1'b1, 1'b0};
1363: data_out = {8'd9, 8'd34, 1'b1, 1'b0};
1364: data_out = {8'd10, 8'd34, 1'b1, 1'b0};
1365: data_out = {8'd11, 8'd34, 1'b1, 1'b0};
1366: data_out = {8'd25, 8'd34, 1'b1, 1'b0};
1367: data_out = {8'd26, 8'd34, 1'b1, 1'b0};
1368: data_out = {8'd27, 8'd34, 1'b1, 1'b0};
1369: data_out = {8'd28, 8'd34, 1'b1, 1'b0};
1370: data_out = {8'd29, 8'd34, 1'b1, 1'b0};
1371: data_out = {8'd30, 8'd34, 1'b1, 1'b0};
1372: data_out = {8'd36, 8'd34, 1'b1, 1'b0};
1373: data_out = {8'd37, 8'd34, 1'b1, 1'b0};
1374: data_out = {8'd38, 8'd34, 1'b1, 1'b0};
1375: data_out = {8'd39, 8'd34, 1'b1, 1'b0};
1376: data_out = {8'd40, 8'd34, 1'b1, 1'b0};
1377: data_out = {8'd41, 8'd34, 1'b1, 1'b0};
1378: data_out = {8'd55, 8'd34, 1'b1, 1'b0};
1379: data_out = {8'd56, 8'd34, 1'b1, 1'b0};
1380: data_out = {8'd57, 8'd34, 1'b1, 1'b0};
1381: data_out = {8'd58, 8'd34, 1'b1, 1'b0};
1382: data_out = {8'd59, 8'd34, 1'b1, 1'b0};
1383: data_out = {8'd60, 8'd34, 1'b1, 1'b0};
1384: data_out = {8'd73, 8'd34, 1'b1, 1'b0};
1385: data_out = {8'd74, 8'd34, 1'b1, 1'b0};
1386: data_out = {8'd75, 8'd34, 1'b1, 1'b0};
1387: data_out = {8'd76, 8'd34, 1'b1, 1'b0};
1388: data_out = {8'd77, 8'd34, 1'b1, 1'b0};
1389: data_out = {8'd78, 8'd34, 1'b1, 1'b0};
1390: data_out = {8'd107, 8'd34, 1'b1, 1'b0};
1391: data_out = {8'd108, 8'd34, 1'b1, 1'b0};
1392: data_out = {8'd109, 8'd34, 1'b1, 1'b0};
1393: data_out = {8'd110, 8'd34, 1'b1, 1'b0};
1394: data_out = {8'd111, 8'd34, 1'b1, 1'b0};
1395: data_out = {8'd112, 8'd34, 1'b1, 1'b0};
1396: data_out = {8'd113, 8'd34, 1'b1, 1'b0};
1397: data_out = {8'd114, 8'd34, 1'b1, 1'b0};
1398: data_out = {8'd115, 8'd34, 1'b1, 1'b0};
1399: data_out = {8'd116, 8'd34, 1'b1, 1'b0};
1400: data_out = {8'd117, 8'd34, 1'b1, 1'b0};
1401: data_out = {8'd118, 8'd34, 1'b1, 1'b0};
1402: data_out = {8'd119, 8'd34, 1'b1, 1'b0};
1403: data_out = {8'd120, 8'd34, 1'b1, 1'b0};
1404: data_out = {8'd121, 8'd34, 1'b1, 1'b0};
1405: data_out = {8'd127, 8'd34, 1'b1, 1'b0};
1406: data_out = {8'd128, 8'd34, 1'b1, 1'b0};
1407: data_out = {8'd129, 8'd34, 1'b1, 1'b0};
1408: data_out = {8'd130, 8'd34, 1'b1, 1'b0};
1409: data_out = {8'd131, 8'd34, 1'b1, 1'b0};
1410: data_out = {8'd132, 8'd34, 1'b1, 1'b0};
1411: data_out = {8'd146, 8'd34, 1'b1, 1'b0};
1412: data_out = {8'd147, 8'd34, 1'b1, 1'b0};
1413: data_out = {8'd148, 8'd34, 1'b1, 1'b0};
1414: data_out = {8'd149, 8'd34, 1'b1, 1'b0};
1415: data_out = {8'd150, 8'd34, 1'b1, 1'b0};
1416: data_out = {8'd151, 8'd34, 1'b1, 1'b0};
1417: data_out = {8'd160, 8'd34, 1'b1, 1'b0};
1418: data_out = {8'd161, 8'd34, 1'b1, 1'b0};
1419: data_out = {8'd162, 8'd34, 1'b1, 1'b0};
1420: data_out = {8'd163, 8'd34, 1'b1, 1'b0};
1421: data_out = {8'd164, 8'd34, 1'b1, 1'b0};
1422: data_out = {8'd165, 8'd34, 1'b1, 1'b0};
1423: data_out = {8'd166, 8'd34, 1'b1, 1'b0};
1424: data_out = {8'd167, 8'd34, 1'b1, 1'b0};
1425: data_out = {8'd168, 8'd34, 1'b1, 1'b0};
1426: data_out = {8'd169, 8'd34, 1'b1, 1'b0};
1427: data_out = {8'd170, 8'd34, 1'b1, 1'b0};
1428: data_out = {8'd171, 8'd34, 1'b1, 1'b0};
1429: data_out = {8'd172, 8'd34, 1'b1, 1'b0};
1430: data_out = {8'd173, 8'd34, 1'b1, 1'b0};
1431: data_out = {8'd174, 8'd34, 1'b1, 1'b0};
1432: data_out = {8'd175, 8'd34, 1'b1, 1'b0};
1433: data_out = {8'd176, 8'd34, 1'b1, 1'b0};
1434: data_out = {8'd177, 8'd34, 1'b1, 1'b0};
1435: data_out = {8'd178, 8'd34, 1'b1, 1'b0};
1436: data_out = {8'd197, 8'd34, 1'b1, 1'b0};
1437: data_out = {8'd198, 8'd34, 1'b1, 1'b0};
1438: data_out = {8'd199, 8'd34, 1'b1, 1'b0};
1439: data_out = {8'd200, 8'd34, 1'b1, 1'b0};
1440: data_out = {8'd201, 8'd34, 1'b1, 1'b0};
1441: data_out = {8'd202, 8'd34, 1'b1, 1'b0};
1442: data_out = {8'd203, 8'd34, 1'b1, 1'b0};
1443: data_out = {8'd204, 8'd34, 1'b1, 1'b0};
1444: data_out = {8'd205, 8'd34, 1'b1, 1'b0};
1445: data_out = {8'd206, 8'd34, 1'b1, 1'b0};
1446: data_out = {8'd207, 8'd34, 1'b1, 1'b0};
1447: data_out = {8'd208, 8'd34, 1'b1, 1'b0};
1448: data_out = {8'd209, 8'd34, 1'b1, 1'b0};
1449: data_out = {8'd210, 8'd34, 1'b1, 1'b0};
1450: data_out = {8'd211, 8'd34, 1'b1, 1'b0};
1451: data_out = {8'd6, 8'd35, 1'b1, 1'b0};
1452: data_out = {8'd7, 8'd35, 1'b1, 1'b0};
1453: data_out = {8'd8, 8'd35, 1'b1, 1'b0};
1454: data_out = {8'd9, 8'd35, 1'b1, 1'b0};
1455: data_out = {8'd10, 8'd35, 1'b1, 1'b0};
1456: data_out = {8'd11, 8'd35, 1'b1, 1'b0};
1457: data_out = {8'd25, 8'd35, 1'b1, 1'b0};
1458: data_out = {8'd26, 8'd35, 1'b1, 1'b0};
1459: data_out = {8'd27, 8'd35, 1'b1, 1'b0};
1460: data_out = {8'd28, 8'd35, 1'b1, 1'b0};
1461: data_out = {8'd29, 8'd35, 1'b1, 1'b0};
1462: data_out = {8'd30, 8'd35, 1'b1, 1'b0};
1463: data_out = {8'd36, 8'd35, 1'b1, 1'b0};
1464: data_out = {8'd37, 8'd35, 1'b1, 1'b0};
1465: data_out = {8'd38, 8'd35, 1'b1, 1'b0};
1466: data_out = {8'd39, 8'd35, 1'b1, 1'b0};
1467: data_out = {8'd40, 8'd35, 1'b1, 1'b0};
1468: data_out = {8'd41, 8'd35, 1'b1, 1'b0};
1469: data_out = {8'd55, 8'd35, 1'b1, 1'b0};
1470: data_out = {8'd56, 8'd35, 1'b1, 1'b0};
1471: data_out = {8'd57, 8'd35, 1'b1, 1'b0};
1472: data_out = {8'd58, 8'd35, 1'b1, 1'b0};
1473: data_out = {8'd59, 8'd35, 1'b1, 1'b0};
1474: data_out = {8'd60, 8'd35, 1'b1, 1'b0};
1475: data_out = {8'd73, 8'd35, 1'b1, 1'b0};
1476: data_out = {8'd74, 8'd35, 1'b1, 1'b0};
1477: data_out = {8'd75, 8'd35, 1'b1, 1'b0};
1478: data_out = {8'd76, 8'd35, 1'b1, 1'b0};
1479: data_out = {8'd77, 8'd35, 1'b1, 1'b0};
1480: data_out = {8'd78, 8'd35, 1'b1, 1'b0};
1481: data_out = {8'd101, 8'd35, 1'b1, 1'b0};
1482: data_out = {8'd102, 8'd35, 1'b1, 1'b0};
1483: data_out = {8'd103, 8'd35, 1'b1, 1'b0};
1484: data_out = {8'd104, 8'd35, 1'b1, 1'b0};
1485: data_out = {8'd105, 8'd35, 1'b1, 1'b0};
1486: data_out = {8'd106, 8'd35, 1'b1, 1'b0};
1487: data_out = {8'd107, 8'd35, 1'b1, 1'b0};
1488: data_out = {8'd108, 8'd35, 1'b1, 1'b0};
1489: data_out = {8'd109, 8'd35, 1'b1, 1'b0};
1490: data_out = {8'd110, 8'd35, 1'b1, 1'b0};
1491: data_out = {8'd111, 8'd35, 1'b1, 1'b0};
1492: data_out = {8'd112, 8'd35, 1'b1, 1'b0};
1493: data_out = {8'd113, 8'd35, 1'b1, 1'b0};
1494: data_out = {8'd114, 8'd35, 1'b1, 1'b0};
1495: data_out = {8'd115, 8'd35, 1'b1, 1'b0};
1496: data_out = {8'd116, 8'd35, 1'b1, 1'b0};
1497: data_out = {8'd117, 8'd35, 1'b1, 1'b0};
1498: data_out = {8'd118, 8'd35, 1'b1, 1'b0};
1499: data_out = {8'd119, 8'd35, 1'b1, 1'b0};
1500: data_out = {8'd120, 8'd35, 1'b1, 1'b0};
1501: data_out = {8'd121, 8'd35, 1'b1, 1'b0};
1502: data_out = {8'd127, 8'd35, 1'b1, 1'b0};
1503: data_out = {8'd128, 8'd35, 1'b1, 1'b0};
1504: data_out = {8'd129, 8'd35, 1'b1, 1'b0};
1505: data_out = {8'd130, 8'd35, 1'b1, 1'b0};
1506: data_out = {8'd131, 8'd35, 1'b1, 1'b0};
1507: data_out = {8'd132, 8'd35, 1'b1, 1'b0};
1508: data_out = {8'd146, 8'd35, 1'b1, 1'b0};
1509: data_out = {8'd147, 8'd35, 1'b1, 1'b0};
1510: data_out = {8'd148, 8'd35, 1'b1, 1'b0};
1511: data_out = {8'd149, 8'd35, 1'b1, 1'b0};
1512: data_out = {8'd150, 8'd35, 1'b1, 1'b0};
1513: data_out = {8'd151, 8'd35, 1'b1, 1'b0};
1514: data_out = {8'd160, 8'd35, 1'b1, 1'b0};
1515: data_out = {8'd161, 8'd35, 1'b1, 1'b0};
1516: data_out = {8'd162, 8'd35, 1'b1, 1'b0};
1517: data_out = {8'd163, 8'd35, 1'b1, 1'b0};
1518: data_out = {8'd164, 8'd35, 1'b1, 1'b0};
1519: data_out = {8'd165, 8'd35, 1'b1, 1'b0};
1520: data_out = {8'd166, 8'd35, 1'b1, 1'b0};
1521: data_out = {8'd167, 8'd35, 1'b1, 1'b0};
1522: data_out = {8'd168, 8'd35, 1'b1, 1'b0};
1523: data_out = {8'd169, 8'd35, 1'b1, 1'b0};
1524: data_out = {8'd170, 8'd35, 1'b1, 1'b0};
1525: data_out = {8'd171, 8'd35, 1'b1, 1'b0};
1526: data_out = {8'd172, 8'd35, 1'b1, 1'b0};
1527: data_out = {8'd173, 8'd35, 1'b1, 1'b0};
1528: data_out = {8'd174, 8'd35, 1'b1, 1'b0};
1529: data_out = {8'd175, 8'd35, 1'b1, 1'b0};
1530: data_out = {8'd176, 8'd35, 1'b1, 1'b0};
1531: data_out = {8'd177, 8'd35, 1'b1, 1'b0};
1532: data_out = {8'd178, 8'd35, 1'b1, 1'b0};
1533: data_out = {8'd191, 8'd35, 1'b1, 1'b0};
1534: data_out = {8'd192, 8'd35, 1'b1, 1'b0};
1535: data_out = {8'd193, 8'd35, 1'b1, 1'b0};
1536: data_out = {8'd194, 8'd35, 1'b1, 1'b0};
1537: data_out = {8'd195, 8'd35, 1'b1, 1'b0};
1538: data_out = {8'd196, 8'd35, 1'b1, 1'b0};
1539: data_out = {8'd197, 8'd35, 1'b1, 1'b0};
1540: data_out = {8'd198, 8'd35, 1'b1, 1'b0};
1541: data_out = {8'd199, 8'd35, 1'b1, 1'b0};
1542: data_out = {8'd200, 8'd35, 1'b1, 1'b0};
1543: data_out = {8'd201, 8'd35, 1'b1, 1'b0};
1544: data_out = {8'd202, 8'd35, 1'b1, 1'b0};
1545: data_out = {8'd203, 8'd35, 1'b1, 1'b0};
1546: data_out = {8'd204, 8'd35, 1'b1, 1'b0};
1547: data_out = {8'd205, 8'd35, 1'b1, 1'b0};
1548: data_out = {8'd206, 8'd35, 1'b1, 1'b0};
1549: data_out = {8'd207, 8'd35, 1'b1, 1'b0};
1550: data_out = {8'd208, 8'd35, 1'b1, 1'b0};
1551: data_out = {8'd209, 8'd35, 1'b1, 1'b0};
1552: data_out = {8'd210, 8'd35, 1'b1, 1'b0};
1553: data_out = {8'd211, 8'd35, 1'b1, 1'b0};
1554: data_out = {8'd6, 8'd36, 1'b1, 1'b0};
1555: data_out = {8'd7, 8'd36, 1'b1, 1'b0};
1556: data_out = {8'd8, 8'd36, 1'b1, 1'b0};
1557: data_out = {8'd9, 8'd36, 1'b1, 1'b0};
1558: data_out = {8'd10, 8'd36, 1'b1, 1'b0};
1559: data_out = {8'd11, 8'd36, 1'b1, 1'b0};
1560: data_out = {8'd25, 8'd36, 1'b1, 1'b0};
1561: data_out = {8'd26, 8'd36, 1'b1, 1'b0};
1562: data_out = {8'd27, 8'd36, 1'b1, 1'b0};
1563: data_out = {8'd28, 8'd36, 1'b1, 1'b0};
1564: data_out = {8'd29, 8'd36, 1'b1, 1'b0};
1565: data_out = {8'd30, 8'd36, 1'b1, 1'b0};
1566: data_out = {8'd36, 8'd36, 1'b1, 1'b0};
1567: data_out = {8'd37, 8'd36, 1'b1, 1'b0};
1568: data_out = {8'd38, 8'd36, 1'b1, 1'b0};
1569: data_out = {8'd39, 8'd36, 1'b1, 1'b0};
1570: data_out = {8'd40, 8'd36, 1'b1, 1'b0};
1571: data_out = {8'd41, 8'd36, 1'b1, 1'b0};
1572: data_out = {8'd55, 8'd36, 1'b1, 1'b0};
1573: data_out = {8'd56, 8'd36, 1'b1, 1'b0};
1574: data_out = {8'd57, 8'd36, 1'b1, 1'b0};
1575: data_out = {8'd58, 8'd36, 1'b1, 1'b0};
1576: data_out = {8'd59, 8'd36, 1'b1, 1'b0};
1577: data_out = {8'd60, 8'd36, 1'b1, 1'b0};
1578: data_out = {8'd73, 8'd36, 1'b1, 1'b0};
1579: data_out = {8'd74, 8'd36, 1'b1, 1'b0};
1580: data_out = {8'd75, 8'd36, 1'b1, 1'b0};
1581: data_out = {8'd76, 8'd36, 1'b1, 1'b0};
1582: data_out = {8'd77, 8'd36, 1'b1, 1'b0};
1583: data_out = {8'd78, 8'd36, 1'b1, 1'b0};
1584: data_out = {8'd98, 8'd36, 1'b1, 1'b0};
1585: data_out = {8'd99, 8'd36, 1'b1, 1'b0};
1586: data_out = {8'd100, 8'd36, 1'b1, 1'b0};
1587: data_out = {8'd101, 8'd36, 1'b1, 1'b0};
1588: data_out = {8'd102, 8'd36, 1'b1, 1'b0};
1589: data_out = {8'd103, 8'd36, 1'b1, 1'b0};
1590: data_out = {8'd104, 8'd36, 1'b1, 1'b0};
1591: data_out = {8'd105, 8'd36, 1'b1, 1'b0};
1592: data_out = {8'd106, 8'd36, 1'b1, 1'b0};
1593: data_out = {8'd107, 8'd36, 1'b1, 1'b0};
1594: data_out = {8'd108, 8'd36, 1'b1, 1'b0};
1595: data_out = {8'd109, 8'd36, 1'b1, 1'b0};
1596: data_out = {8'd110, 8'd36, 1'b1, 1'b0};
1597: data_out = {8'd111, 8'd36, 1'b1, 1'b0};
1598: data_out = {8'd112, 8'd36, 1'b1, 1'b0};
1599: data_out = {8'd113, 8'd36, 1'b1, 1'b0};
1600: data_out = {8'd114, 8'd36, 1'b1, 1'b0};
1601: data_out = {8'd115, 8'd36, 1'b1, 1'b0};
1602: data_out = {8'd116, 8'd36, 1'b1, 1'b0};
1603: data_out = {8'd117, 8'd36, 1'b1, 1'b0};
1604: data_out = {8'd118, 8'd36, 1'b1, 1'b0};
1605: data_out = {8'd119, 8'd36, 1'b1, 1'b0};
1606: data_out = {8'd120, 8'd36, 1'b1, 1'b0};
1607: data_out = {8'd121, 8'd36, 1'b1, 1'b0};
1608: data_out = {8'd127, 8'd36, 1'b1, 1'b0};
1609: data_out = {8'd128, 8'd36, 1'b1, 1'b0};
1610: data_out = {8'd129, 8'd36, 1'b1, 1'b0};
1611: data_out = {8'd130, 8'd36, 1'b1, 1'b0};
1612: data_out = {8'd131, 8'd36, 1'b1, 1'b0};
1613: data_out = {8'd132, 8'd36, 1'b1, 1'b0};
1614: data_out = {8'd146, 8'd36, 1'b1, 1'b0};
1615: data_out = {8'd147, 8'd36, 1'b1, 1'b0};
1616: data_out = {8'd148, 8'd36, 1'b1, 1'b0};
1617: data_out = {8'd149, 8'd36, 1'b1, 1'b0};
1618: data_out = {8'd150, 8'd36, 1'b1, 1'b0};
1619: data_out = {8'd151, 8'd36, 1'b1, 1'b0};
1620: data_out = {8'd160, 8'd36, 1'b1, 1'b0};
1621: data_out = {8'd161, 8'd36, 1'b1, 1'b0};
1622: data_out = {8'd162, 8'd36, 1'b1, 1'b0};
1623: data_out = {8'd163, 8'd36, 1'b1, 1'b0};
1624: data_out = {8'd164, 8'd36, 1'b1, 1'b0};
1625: data_out = {8'd165, 8'd36, 1'b1, 1'b0};
1626: data_out = {8'd166, 8'd36, 1'b1, 1'b0};
1627: data_out = {8'd167, 8'd36, 1'b1, 1'b0};
1628: data_out = {8'd168, 8'd36, 1'b1, 1'b0};
1629: data_out = {8'd169, 8'd36, 1'b1, 1'b0};
1630: data_out = {8'd170, 8'd36, 1'b1, 1'b0};
1631: data_out = {8'd171, 8'd36, 1'b1, 1'b0};
1632: data_out = {8'd172, 8'd36, 1'b1, 1'b0};
1633: data_out = {8'd173, 8'd36, 1'b1, 1'b0};
1634: data_out = {8'd174, 8'd36, 1'b1, 1'b0};
1635: data_out = {8'd175, 8'd36, 1'b1, 1'b0};
1636: data_out = {8'd176, 8'd36, 1'b1, 1'b0};
1637: data_out = {8'd177, 8'd36, 1'b1, 1'b0};
1638: data_out = {8'd178, 8'd36, 1'b1, 1'b0};
1639: data_out = {8'd188, 8'd36, 1'b1, 1'b0};
1640: data_out = {8'd189, 8'd36, 1'b1, 1'b0};
1641: data_out = {8'd190, 8'd36, 1'b1, 1'b0};
1642: data_out = {8'd191, 8'd36, 1'b1, 1'b0};
1643: data_out = {8'd192, 8'd36, 1'b1, 1'b0};
1644: data_out = {8'd193, 8'd36, 1'b1, 1'b0};
1645: data_out = {8'd194, 8'd36, 1'b1, 1'b0};
1646: data_out = {8'd195, 8'd36, 1'b1, 1'b0};
1647: data_out = {8'd196, 8'd36, 1'b1, 1'b0};
1648: data_out = {8'd197, 8'd36, 1'b1, 1'b0};
1649: data_out = {8'd198, 8'd36, 1'b1, 1'b0};
1650: data_out = {8'd199, 8'd36, 1'b1, 1'b0};
1651: data_out = {8'd200, 8'd36, 1'b1, 1'b0};
1652: data_out = {8'd201, 8'd36, 1'b1, 1'b0};
1653: data_out = {8'd202, 8'd36, 1'b1, 1'b0};
1654: data_out = {8'd203, 8'd36, 1'b1, 1'b0};
1655: data_out = {8'd204, 8'd36, 1'b1, 1'b0};
1656: data_out = {8'd205, 8'd36, 1'b1, 1'b0};
1657: data_out = {8'd206, 8'd36, 1'b1, 1'b0};
1658: data_out = {8'd207, 8'd36, 1'b1, 1'b0};
1659: data_out = {8'd208, 8'd36, 1'b1, 1'b0};
1660: data_out = {8'd209, 8'd36, 1'b1, 1'b0};
1661: data_out = {8'd210, 8'd36, 1'b1, 1'b0};
1662: data_out = {8'd211, 8'd36, 1'b1, 1'b0};
1663: data_out = {8'd6, 8'd37, 1'b1, 1'b0};
1664: data_out = {8'd7, 8'd37, 1'b1, 1'b0};
1665: data_out = {8'd8, 8'd37, 1'b1, 1'b0};
1666: data_out = {8'd9, 8'd37, 1'b1, 1'b0};
1667: data_out = {8'd10, 8'd37, 1'b1, 1'b0};
1668: data_out = {8'd11, 8'd37, 1'b1, 1'b0};
1669: data_out = {8'd25, 8'd37, 1'b1, 1'b0};
1670: data_out = {8'd26, 8'd37, 1'b1, 1'b0};
1671: data_out = {8'd27, 8'd37, 1'b1, 1'b0};
1672: data_out = {8'd28, 8'd37, 1'b1, 1'b0};
1673: data_out = {8'd29, 8'd37, 1'b1, 1'b0};
1674: data_out = {8'd30, 8'd37, 1'b1, 1'b0};
1675: data_out = {8'd36, 8'd37, 1'b1, 1'b0};
1676: data_out = {8'd37, 8'd37, 1'b1, 1'b0};
1677: data_out = {8'd38, 8'd37, 1'b1, 1'b0};
1678: data_out = {8'd39, 8'd37, 1'b1, 1'b0};
1679: data_out = {8'd40, 8'd37, 1'b1, 1'b0};
1680: data_out = {8'd41, 8'd37, 1'b1, 1'b0};
1681: data_out = {8'd55, 8'd37, 1'b1, 1'b0};
1682: data_out = {8'd56, 8'd37, 1'b1, 1'b0};
1683: data_out = {8'd57, 8'd37, 1'b1, 1'b0};
1684: data_out = {8'd58, 8'd37, 1'b1, 1'b0};
1685: data_out = {8'd59, 8'd37, 1'b1, 1'b0};
1686: data_out = {8'd60, 8'd37, 1'b1, 1'b0};
1687: data_out = {8'd73, 8'd37, 1'b1, 1'b0};
1688: data_out = {8'd74, 8'd37, 1'b1, 1'b0};
1689: data_out = {8'd75, 8'd37, 1'b1, 1'b0};
1690: data_out = {8'd76, 8'd37, 1'b1, 1'b0};
1691: data_out = {8'd77, 8'd37, 1'b1, 1'b0};
1692: data_out = {8'd78, 8'd37, 1'b1, 1'b0};
1693: data_out = {8'd97, 8'd37, 1'b1, 1'b0};
1694: data_out = {8'd98, 8'd37, 1'b1, 1'b0};
1695: data_out = {8'd99, 8'd37, 1'b1, 1'b0};
1696: data_out = {8'd100, 8'd37, 1'b1, 1'b0};
1697: data_out = {8'd101, 8'd37, 1'b1, 1'b0};
1698: data_out = {8'd102, 8'd37, 1'b1, 1'b0};
1699: data_out = {8'd103, 8'd37, 1'b1, 1'b0};
1700: data_out = {8'd104, 8'd37, 1'b1, 1'b0};
1701: data_out = {8'd105, 8'd37, 1'b1, 1'b0};
1702: data_out = {8'd106, 8'd37, 1'b1, 1'b0};
1703: data_out = {8'd107, 8'd37, 1'b1, 1'b0};
1704: data_out = {8'd108, 8'd37, 1'b1, 1'b0};
1705: data_out = {8'd109, 8'd37, 1'b1, 1'b0};
1706: data_out = {8'd110, 8'd37, 1'b1, 1'b0};
1707: data_out = {8'd111, 8'd37, 1'b1, 1'b0};
1708: data_out = {8'd112, 8'd37, 1'b1, 1'b0};
1709: data_out = {8'd113, 8'd37, 1'b1, 1'b0};
1710: data_out = {8'd114, 8'd37, 1'b1, 1'b0};
1711: data_out = {8'd115, 8'd37, 1'b1, 1'b0};
1712: data_out = {8'd116, 8'd37, 1'b1, 1'b0};
1713: data_out = {8'd117, 8'd37, 1'b1, 1'b0};
1714: data_out = {8'd118, 8'd37, 1'b1, 1'b0};
1715: data_out = {8'd119, 8'd37, 1'b1, 1'b0};
1716: data_out = {8'd120, 8'd37, 1'b1, 1'b0};
1717: data_out = {8'd121, 8'd37, 1'b1, 1'b0};
1718: data_out = {8'd127, 8'd37, 1'b1, 1'b0};
1719: data_out = {8'd128, 8'd37, 1'b1, 1'b0};
1720: data_out = {8'd129, 8'd37, 1'b1, 1'b0};
1721: data_out = {8'd130, 8'd37, 1'b1, 1'b0};
1722: data_out = {8'd131, 8'd37, 1'b1, 1'b0};
1723: data_out = {8'd132, 8'd37, 1'b1, 1'b0};
1724: data_out = {8'd146, 8'd37, 1'b1, 1'b0};
1725: data_out = {8'd147, 8'd37, 1'b1, 1'b0};
1726: data_out = {8'd148, 8'd37, 1'b1, 1'b0};
1727: data_out = {8'd149, 8'd37, 1'b1, 1'b0};
1728: data_out = {8'd150, 8'd37, 1'b1, 1'b0};
1729: data_out = {8'd151, 8'd37, 1'b1, 1'b0};
1730: data_out = {8'd160, 8'd37, 1'b1, 1'b0};
1731: data_out = {8'd161, 8'd37, 1'b1, 1'b0};
1732: data_out = {8'd162, 8'd37, 1'b1, 1'b0};
1733: data_out = {8'd163, 8'd37, 1'b1, 1'b0};
1734: data_out = {8'd164, 8'd37, 1'b1, 1'b0};
1735: data_out = {8'd165, 8'd37, 1'b1, 1'b0};
1736: data_out = {8'd166, 8'd37, 1'b1, 1'b0};
1737: data_out = {8'd167, 8'd37, 1'b1, 1'b0};
1738: data_out = {8'd168, 8'd37, 1'b1, 1'b0};
1739: data_out = {8'd169, 8'd37, 1'b1, 1'b0};
1740: data_out = {8'd170, 8'd37, 1'b1, 1'b0};
1741: data_out = {8'd171, 8'd37, 1'b1, 1'b0};
1742: data_out = {8'd172, 8'd37, 1'b1, 1'b0};
1743: data_out = {8'd173, 8'd37, 1'b1, 1'b0};
1744: data_out = {8'd174, 8'd37, 1'b1, 1'b0};
1745: data_out = {8'd175, 8'd37, 1'b1, 1'b0};
1746: data_out = {8'd176, 8'd37, 1'b1, 1'b0};
1747: data_out = {8'd177, 8'd37, 1'b1, 1'b0};
1748: data_out = {8'd178, 8'd37, 1'b1, 1'b0};
1749: data_out = {8'd187, 8'd37, 1'b1, 1'b0};
1750: data_out = {8'd188, 8'd37, 1'b1, 1'b0};
1751: data_out = {8'd189, 8'd37, 1'b1, 1'b0};
1752: data_out = {8'd190, 8'd37, 1'b1, 1'b0};
1753: data_out = {8'd191, 8'd37, 1'b1, 1'b0};
1754: data_out = {8'd192, 8'd37, 1'b1, 1'b0};
1755: data_out = {8'd193, 8'd37, 1'b1, 1'b0};
1756: data_out = {8'd194, 8'd37, 1'b1, 1'b0};
1757: data_out = {8'd195, 8'd37, 1'b1, 1'b0};
1758: data_out = {8'd196, 8'd37, 1'b1, 1'b0};
1759: data_out = {8'd197, 8'd37, 1'b1, 1'b0};
1760: data_out = {8'd198, 8'd37, 1'b1, 1'b0};
1761: data_out = {8'd199, 8'd37, 1'b1, 1'b0};
1762: data_out = {8'd200, 8'd37, 1'b1, 1'b0};
1763: data_out = {8'd201, 8'd37, 1'b1, 1'b0};
1764: data_out = {8'd202, 8'd37, 1'b1, 1'b0};
1765: data_out = {8'd203, 8'd37, 1'b1, 1'b0};
1766: data_out = {8'd204, 8'd37, 1'b1, 1'b0};
1767: data_out = {8'd205, 8'd37, 1'b1, 1'b0};
1768: data_out = {8'd206, 8'd37, 1'b1, 1'b0};
1769: data_out = {8'd207, 8'd37, 1'b1, 1'b0};
1770: data_out = {8'd208, 8'd37, 1'b1, 1'b0};
1771: data_out = {8'd209, 8'd37, 1'b1, 1'b0};
1772: data_out = {8'd210, 8'd37, 1'b1, 1'b0};
1773: data_out = {8'd211, 8'd37, 1'b1, 1'b0};
1774: data_out = {8'd6, 8'd38, 1'b1, 1'b0};
1775: data_out = {8'd7, 8'd38, 1'b1, 1'b0};
1776: data_out = {8'd8, 8'd38, 1'b1, 1'b0};
1777: data_out = {8'd9, 8'd38, 1'b1, 1'b0};
1778: data_out = {8'd10, 8'd38, 1'b1, 1'b0};
1779: data_out = {8'd11, 8'd38, 1'b1, 1'b0};
1780: data_out = {8'd25, 8'd38, 1'b1, 1'b0};
1781: data_out = {8'd26, 8'd38, 1'b1, 1'b0};
1782: data_out = {8'd27, 8'd38, 1'b1, 1'b0};
1783: data_out = {8'd28, 8'd38, 1'b1, 1'b0};
1784: data_out = {8'd29, 8'd38, 1'b1, 1'b0};
1785: data_out = {8'd30, 8'd38, 1'b1, 1'b0};
1786: data_out = {8'd36, 8'd38, 1'b1, 1'b0};
1787: data_out = {8'd37, 8'd38, 1'b1, 1'b0};
1788: data_out = {8'd38, 8'd38, 1'b1, 1'b0};
1789: data_out = {8'd39, 8'd38, 1'b1, 1'b0};
1790: data_out = {8'd40, 8'd38, 1'b1, 1'b0};
1791: data_out = {8'd41, 8'd38, 1'b1, 1'b0};
1792: data_out = {8'd55, 8'd38, 1'b1, 1'b0};
1793: data_out = {8'd56, 8'd38, 1'b1, 1'b0};
1794: data_out = {8'd57, 8'd38, 1'b1, 1'b0};
1795: data_out = {8'd58, 8'd38, 1'b1, 1'b0};
1796: data_out = {8'd59, 8'd38, 1'b1, 1'b0};
1797: data_out = {8'd60, 8'd38, 1'b1, 1'b0};
1798: data_out = {8'd73, 8'd38, 1'b1, 1'b0};
1799: data_out = {8'd74, 8'd38, 1'b1, 1'b0};
1800: data_out = {8'd75, 8'd38, 1'b1, 1'b0};
1801: data_out = {8'd76, 8'd38, 1'b1, 1'b0};
1802: data_out = {8'd77, 8'd38, 1'b1, 1'b0};
1803: data_out = {8'd78, 8'd38, 1'b1, 1'b0};
1804: data_out = {8'd97, 8'd38, 1'b1, 1'b0};
1805: data_out = {8'd98, 8'd38, 1'b1, 1'b0};
1806: data_out = {8'd99, 8'd38, 1'b1, 1'b0};
1807: data_out = {8'd100, 8'd38, 1'b1, 1'b0};
1808: data_out = {8'd101, 8'd38, 1'b1, 1'b0};
1809: data_out = {8'd102, 8'd38, 1'b1, 1'b0};
1810: data_out = {8'd103, 8'd38, 1'b1, 1'b0};
1811: data_out = {8'd104, 8'd38, 1'b1, 1'b0};
1812: data_out = {8'd105, 8'd38, 1'b1, 1'b0};
1813: data_out = {8'd106, 8'd38, 1'b1, 1'b0};
1814: data_out = {8'd107, 8'd38, 1'b1, 1'b0};
1815: data_out = {8'd108, 8'd38, 1'b1, 1'b0};
1816: data_out = {8'd109, 8'd38, 1'b1, 1'b0};
1817: data_out = {8'd116, 8'd38, 1'b1, 1'b0};
1818: data_out = {8'd117, 8'd38, 1'b1, 1'b0};
1819: data_out = {8'd118, 8'd38, 1'b1, 1'b0};
1820: data_out = {8'd119, 8'd38, 1'b1, 1'b0};
1821: data_out = {8'd120, 8'd38, 1'b1, 1'b0};
1822: data_out = {8'd121, 8'd38, 1'b1, 1'b0};
1823: data_out = {8'd127, 8'd38, 1'b1, 1'b0};
1824: data_out = {8'd128, 8'd38, 1'b1, 1'b0};
1825: data_out = {8'd129, 8'd38, 1'b1, 1'b0};
1826: data_out = {8'd130, 8'd38, 1'b1, 1'b0};
1827: data_out = {8'd131, 8'd38, 1'b1, 1'b0};
1828: data_out = {8'd132, 8'd38, 1'b1, 1'b0};
1829: data_out = {8'd146, 8'd38, 1'b1, 1'b0};
1830: data_out = {8'd147, 8'd38, 1'b1, 1'b0};
1831: data_out = {8'd148, 8'd38, 1'b1, 1'b0};
1832: data_out = {8'd149, 8'd38, 1'b1, 1'b0};
1833: data_out = {8'd150, 8'd38, 1'b1, 1'b0};
1834: data_out = {8'd151, 8'd38, 1'b1, 1'b0};
1835: data_out = {8'd160, 8'd38, 1'b1, 1'b0};
1836: data_out = {8'd161, 8'd38, 1'b1, 1'b0};
1837: data_out = {8'd162, 8'd38, 1'b1, 1'b0};
1838: data_out = {8'd163, 8'd38, 1'b1, 1'b0};
1839: data_out = {8'd164, 8'd38, 1'b1, 1'b0};
1840: data_out = {8'd165, 8'd38, 1'b1, 1'b0};
1841: data_out = {8'd166, 8'd38, 1'b1, 1'b0};
1842: data_out = {8'd167, 8'd38, 1'b1, 1'b0};
1843: data_out = {8'd168, 8'd38, 1'b1, 1'b0};
1844: data_out = {8'd169, 8'd38, 1'b1, 1'b0};
1845: data_out = {8'd170, 8'd38, 1'b1, 1'b0};
1846: data_out = {8'd171, 8'd38, 1'b1, 1'b0};
1847: data_out = {8'd172, 8'd38, 1'b1, 1'b0};
1848: data_out = {8'd173, 8'd38, 1'b1, 1'b0};
1849: data_out = {8'd174, 8'd38, 1'b1, 1'b0};
1850: data_out = {8'd175, 8'd38, 1'b1, 1'b0};
1851: data_out = {8'd176, 8'd38, 1'b1, 1'b0};
1852: data_out = {8'd177, 8'd38, 1'b1, 1'b0};
1853: data_out = {8'd178, 8'd38, 1'b1, 1'b0};
1854: data_out = {8'd187, 8'd38, 1'b1, 1'b0};
1855: data_out = {8'd188, 8'd38, 1'b1, 1'b0};
1856: data_out = {8'd189, 8'd38, 1'b1, 1'b0};
1857: data_out = {8'd190, 8'd38, 1'b1, 1'b0};
1858: data_out = {8'd191, 8'd38, 1'b1, 1'b0};
1859: data_out = {8'd192, 8'd38, 1'b1, 1'b0};
1860: data_out = {8'd193, 8'd38, 1'b1, 1'b0};
1861: data_out = {8'd194, 8'd38, 1'b1, 1'b0};
1862: data_out = {8'd195, 8'd38, 1'b1, 1'b0};
1863: data_out = {8'd196, 8'd38, 1'b1, 1'b0};
1864: data_out = {8'd197, 8'd38, 1'b1, 1'b0};
1865: data_out = {8'd198, 8'd38, 1'b1, 1'b0};
1866: data_out = {8'd199, 8'd38, 1'b1, 1'b0};
1867: data_out = {8'd206, 8'd38, 1'b1, 1'b0};
1868: data_out = {8'd207, 8'd38, 1'b1, 1'b0};
1869: data_out = {8'd208, 8'd38, 1'b1, 1'b0};
1870: data_out = {8'd209, 8'd38, 1'b1, 1'b0};
1871: data_out = {8'd210, 8'd38, 1'b1, 1'b0};
1872: data_out = {8'd211, 8'd38, 1'b1, 1'b0};
1873: data_out = {8'd6, 8'd39, 1'b1, 1'b0};
1874: data_out = {8'd7, 8'd39, 1'b1, 1'b0};
1875: data_out = {8'd8, 8'd39, 1'b1, 1'b0};
1876: data_out = {8'd9, 8'd39, 1'b1, 1'b0};
1877: data_out = {8'd10, 8'd39, 1'b1, 1'b0};
1878: data_out = {8'd11, 8'd39, 1'b1, 1'b0};
1879: data_out = {8'd25, 8'd39, 1'b1, 1'b0};
1880: data_out = {8'd26, 8'd39, 1'b1, 1'b0};
1881: data_out = {8'd27, 8'd39, 1'b1, 1'b0};
1882: data_out = {8'd28, 8'd39, 1'b1, 1'b0};
1883: data_out = {8'd29, 8'd39, 1'b1, 1'b0};
1884: data_out = {8'd30, 8'd39, 1'b1, 1'b0};
1885: data_out = {8'd36, 8'd39, 1'b1, 1'b0};
1886: data_out = {8'd37, 8'd39, 1'b1, 1'b0};
1887: data_out = {8'd38, 8'd39, 1'b1, 1'b0};
1888: data_out = {8'd39, 8'd39, 1'b1, 1'b0};
1889: data_out = {8'd40, 8'd39, 1'b1, 1'b0};
1890: data_out = {8'd41, 8'd39, 1'b1, 1'b0};
1891: data_out = {8'd55, 8'd39, 1'b1, 1'b0};
1892: data_out = {8'd56, 8'd39, 1'b1, 1'b0};
1893: data_out = {8'd57, 8'd39, 1'b1, 1'b0};
1894: data_out = {8'd58, 8'd39, 1'b1, 1'b0};
1895: data_out = {8'd59, 8'd39, 1'b1, 1'b0};
1896: data_out = {8'd60, 8'd39, 1'b1, 1'b0};
1897: data_out = {8'd73, 8'd39, 1'b1, 1'b0};
1898: data_out = {8'd74, 8'd39, 1'b1, 1'b0};
1899: data_out = {8'd75, 8'd39, 1'b1, 1'b0};
1900: data_out = {8'd76, 8'd39, 1'b1, 1'b0};
1901: data_out = {8'd77, 8'd39, 1'b1, 1'b0};
1902: data_out = {8'd78, 8'd39, 1'b1, 1'b0};
1903: data_out = {8'd97, 8'd39, 1'b1, 1'b0};
1904: data_out = {8'd98, 8'd39, 1'b1, 1'b0};
1905: data_out = {8'd99, 8'd39, 1'b1, 1'b0};
1906: data_out = {8'd100, 8'd39, 1'b1, 1'b0};
1907: data_out = {8'd101, 8'd39, 1'b1, 1'b0};
1908: data_out = {8'd102, 8'd39, 1'b1, 1'b0};
1909: data_out = {8'd103, 8'd39, 1'b1, 1'b0};
1910: data_out = {8'd104, 8'd39, 1'b1, 1'b0};
1911: data_out = {8'd116, 8'd39, 1'b1, 1'b0};
1912: data_out = {8'd117, 8'd39, 1'b1, 1'b0};
1913: data_out = {8'd118, 8'd39, 1'b1, 1'b0};
1914: data_out = {8'd119, 8'd39, 1'b1, 1'b0};
1915: data_out = {8'd120, 8'd39, 1'b1, 1'b0};
1916: data_out = {8'd121, 8'd39, 1'b1, 1'b0};
1917: data_out = {8'd127, 8'd39, 1'b1, 1'b0};
1918: data_out = {8'd128, 8'd39, 1'b1, 1'b0};
1919: data_out = {8'd129, 8'd39, 1'b1, 1'b0};
1920: data_out = {8'd130, 8'd39, 1'b1, 1'b0};
1921: data_out = {8'd131, 8'd39, 1'b1, 1'b0};
1922: data_out = {8'd132, 8'd39, 1'b1, 1'b0};
1923: data_out = {8'd146, 8'd39, 1'b1, 1'b0};
1924: data_out = {8'd147, 8'd39, 1'b1, 1'b0};
1925: data_out = {8'd148, 8'd39, 1'b1, 1'b0};
1926: data_out = {8'd149, 8'd39, 1'b1, 1'b0};
1927: data_out = {8'd150, 8'd39, 1'b1, 1'b0};
1928: data_out = {8'd151, 8'd39, 1'b1, 1'b0};
1929: data_out = {8'd187, 8'd39, 1'b1, 1'b0};
1930: data_out = {8'd188, 8'd39, 1'b1, 1'b0};
1931: data_out = {8'd189, 8'd39, 1'b1, 1'b0};
1932: data_out = {8'd190, 8'd39, 1'b1, 1'b0};
1933: data_out = {8'd191, 8'd39, 1'b1, 1'b0};
1934: data_out = {8'd192, 8'd39, 1'b1, 1'b0};
1935: data_out = {8'd193, 8'd39, 1'b1, 1'b0};
1936: data_out = {8'd194, 8'd39, 1'b1, 1'b0};
1937: data_out = {8'd206, 8'd39, 1'b1, 1'b0};
1938: data_out = {8'd207, 8'd39, 1'b1, 1'b0};
1939: data_out = {8'd208, 8'd39, 1'b1, 1'b0};
1940: data_out = {8'd209, 8'd39, 1'b1, 1'b0};
1941: data_out = {8'd210, 8'd39, 1'b1, 1'b0};
1942: data_out = {8'd211, 8'd39, 1'b1, 1'b0};
1943: data_out = {8'd6, 8'd40, 1'b1, 1'b0};
1944: data_out = {8'd7, 8'd40, 1'b1, 1'b0};
1945: data_out = {8'd8, 8'd40, 1'b1, 1'b0};
1946: data_out = {8'd9, 8'd40, 1'b1, 1'b0};
1947: data_out = {8'd10, 8'd40, 1'b1, 1'b0};
1948: data_out = {8'd11, 8'd40, 1'b1, 1'b0};
1949: data_out = {8'd25, 8'd40, 1'b1, 1'b0};
1950: data_out = {8'd26, 8'd40, 1'b1, 1'b0};
1951: data_out = {8'd27, 8'd40, 1'b1, 1'b0};
1952: data_out = {8'd28, 8'd40, 1'b1, 1'b0};
1953: data_out = {8'd29, 8'd40, 1'b1, 1'b0};
1954: data_out = {8'd30, 8'd40, 1'b1, 1'b0};
1955: data_out = {8'd36, 8'd40, 1'b1, 1'b0};
1956: data_out = {8'd37, 8'd40, 1'b1, 1'b0};
1957: data_out = {8'd38, 8'd40, 1'b1, 1'b0};
1958: data_out = {8'd39, 8'd40, 1'b1, 1'b0};
1959: data_out = {8'd40, 8'd40, 1'b1, 1'b0};
1960: data_out = {8'd41, 8'd40, 1'b1, 1'b0};
1961: data_out = {8'd55, 8'd40, 1'b1, 1'b0};
1962: data_out = {8'd56, 8'd40, 1'b1, 1'b0};
1963: data_out = {8'd57, 8'd40, 1'b1, 1'b0};
1964: data_out = {8'd58, 8'd40, 1'b1, 1'b0};
1965: data_out = {8'd59, 8'd40, 1'b1, 1'b0};
1966: data_out = {8'd60, 8'd40, 1'b1, 1'b0};
1967: data_out = {8'd73, 8'd40, 1'b1, 1'b0};
1968: data_out = {8'd74, 8'd40, 1'b1, 1'b0};
1969: data_out = {8'd75, 8'd40, 1'b1, 1'b0};
1970: data_out = {8'd76, 8'd40, 1'b1, 1'b0};
1971: data_out = {8'd77, 8'd40, 1'b1, 1'b0};
1972: data_out = {8'd78, 8'd40, 1'b1, 1'b0};
1973: data_out = {8'd97, 8'd40, 1'b1, 1'b0};
1974: data_out = {8'd98, 8'd40, 1'b1, 1'b0};
1975: data_out = {8'd99, 8'd40, 1'b1, 1'b0};
1976: data_out = {8'd100, 8'd40, 1'b1, 1'b0};
1977: data_out = {8'd101, 8'd40, 1'b1, 1'b0};
1978: data_out = {8'd102, 8'd40, 1'b1, 1'b0};
1979: data_out = {8'd116, 8'd40, 1'b1, 1'b0};
1980: data_out = {8'd117, 8'd40, 1'b1, 1'b0};
1981: data_out = {8'd118, 8'd40, 1'b1, 1'b0};
1982: data_out = {8'd119, 8'd40, 1'b1, 1'b0};
1983: data_out = {8'd120, 8'd40, 1'b1, 1'b0};
1984: data_out = {8'd121, 8'd40, 1'b1, 1'b0};
1985: data_out = {8'd127, 8'd40, 1'b1, 1'b0};
1986: data_out = {8'd128, 8'd40, 1'b1, 1'b0};
1987: data_out = {8'd129, 8'd40, 1'b1, 1'b0};
1988: data_out = {8'd130, 8'd40, 1'b1, 1'b0};
1989: data_out = {8'd131, 8'd40, 1'b1, 1'b0};
1990: data_out = {8'd132, 8'd40, 1'b1, 1'b0};
1991: data_out = {8'd146, 8'd40, 1'b1, 1'b0};
1992: data_out = {8'd147, 8'd40, 1'b1, 1'b0};
1993: data_out = {8'd148, 8'd40, 1'b1, 1'b0};
1994: data_out = {8'd149, 8'd40, 1'b1, 1'b0};
1995: data_out = {8'd150, 8'd40, 1'b1, 1'b0};
1996: data_out = {8'd151, 8'd40, 1'b1, 1'b0};
1997: data_out = {8'd187, 8'd40, 1'b1, 1'b0};
1998: data_out = {8'd188, 8'd40, 1'b1, 1'b0};
1999: data_out = {8'd189, 8'd40, 1'b1, 1'b0};
2000: data_out = {8'd190, 8'd40, 1'b1, 1'b0};
2001: data_out = {8'd191, 8'd40, 1'b1, 1'b0};
2002: data_out = {8'd192, 8'd40, 1'b1, 1'b0};
2003: data_out = {8'd206, 8'd40, 1'b1, 1'b0};
2004: data_out = {8'd207, 8'd40, 1'b1, 1'b0};
2005: data_out = {8'd208, 8'd40, 1'b1, 1'b0};
2006: data_out = {8'd209, 8'd40, 1'b1, 1'b0};
2007: data_out = {8'd210, 8'd40, 1'b1, 1'b0};
2008: data_out = {8'd211, 8'd40, 1'b1, 1'b0};
2009: data_out = {8'd6, 8'd41, 1'b1, 1'b0};
2010: data_out = {8'd7, 8'd41, 1'b1, 1'b0};
2011: data_out = {8'd8, 8'd41, 1'b1, 1'b0};
2012: data_out = {8'd9, 8'd41, 1'b1, 1'b0};
2013: data_out = {8'd10, 8'd41, 1'b1, 1'b0};
2014: data_out = {8'd11, 8'd41, 1'b1, 1'b0};
2015: data_out = {8'd25, 8'd41, 1'b1, 1'b0};
2016: data_out = {8'd26, 8'd41, 1'b1, 1'b0};
2017: data_out = {8'd27, 8'd41, 1'b1, 1'b0};
2018: data_out = {8'd28, 8'd41, 1'b1, 1'b0};
2019: data_out = {8'd29, 8'd41, 1'b1, 1'b0};
2020: data_out = {8'd30, 8'd41, 1'b1, 1'b0};
2021: data_out = {8'd36, 8'd41, 1'b1, 1'b0};
2022: data_out = {8'd37, 8'd41, 1'b1, 1'b0};
2023: data_out = {8'd38, 8'd41, 1'b1, 1'b0};
2024: data_out = {8'd39, 8'd41, 1'b1, 1'b0};
2025: data_out = {8'd40, 8'd41, 1'b1, 1'b0};
2026: data_out = {8'd41, 8'd41, 1'b1, 1'b0};
2027: data_out = {8'd55, 8'd41, 1'b1, 1'b0};
2028: data_out = {8'd56, 8'd41, 1'b1, 1'b0};
2029: data_out = {8'd57, 8'd41, 1'b1, 1'b0};
2030: data_out = {8'd58, 8'd41, 1'b1, 1'b0};
2031: data_out = {8'd59, 8'd41, 1'b1, 1'b0};
2032: data_out = {8'd60, 8'd41, 1'b1, 1'b0};
2033: data_out = {8'd73, 8'd41, 1'b1, 1'b0};
2034: data_out = {8'd74, 8'd41, 1'b1, 1'b0};
2035: data_out = {8'd75, 8'd41, 1'b1, 1'b0};
2036: data_out = {8'd76, 8'd41, 1'b1, 1'b0};
2037: data_out = {8'd77, 8'd41, 1'b1, 1'b0};
2038: data_out = {8'd78, 8'd41, 1'b1, 1'b0};
2039: data_out = {8'd97, 8'd41, 1'b1, 1'b0};
2040: data_out = {8'd98, 8'd41, 1'b1, 1'b0};
2041: data_out = {8'd99, 8'd41, 1'b1, 1'b0};
2042: data_out = {8'd100, 8'd41, 1'b1, 1'b0};
2043: data_out = {8'd101, 8'd41, 1'b1, 1'b0};
2044: data_out = {8'd102, 8'd41, 1'b1, 1'b0};
2045: data_out = {8'd116, 8'd41, 1'b1, 1'b0};
2046: data_out = {8'd117, 8'd41, 1'b1, 1'b0};
2047: data_out = {8'd118, 8'd41, 1'b1, 1'b0};
2048: data_out = {8'd119, 8'd41, 1'b1, 1'b0};
2049: data_out = {8'd120, 8'd41, 1'b1, 1'b0};
2050: data_out = {8'd121, 8'd41, 1'b1, 1'b0};
2051: data_out = {8'd127, 8'd41, 1'b1, 1'b0};
2052: data_out = {8'd128, 8'd41, 1'b1, 1'b0};
2053: data_out = {8'd129, 8'd41, 1'b1, 1'b0};
2054: data_out = {8'd130, 8'd41, 1'b1, 1'b0};
2055: data_out = {8'd131, 8'd41, 1'b1, 1'b0};
2056: data_out = {8'd132, 8'd41, 1'b1, 1'b0};
2057: data_out = {8'd146, 8'd41, 1'b1, 1'b0};
2058: data_out = {8'd147, 8'd41, 1'b1, 1'b0};
2059: data_out = {8'd148, 8'd41, 1'b1, 1'b0};
2060: data_out = {8'd149, 8'd41, 1'b1, 1'b0};
2061: data_out = {8'd150, 8'd41, 1'b1, 1'b0};
2062: data_out = {8'd151, 8'd41, 1'b1, 1'b0};
2063: data_out = {8'd187, 8'd41, 1'b1, 1'b0};
2064: data_out = {8'd188, 8'd41, 1'b1, 1'b0};
2065: data_out = {8'd189, 8'd41, 1'b1, 1'b0};
2066: data_out = {8'd190, 8'd41, 1'b1, 1'b0};
2067: data_out = {8'd191, 8'd41, 1'b1, 1'b0};
2068: data_out = {8'd192, 8'd41, 1'b1, 1'b0};
2069: data_out = {8'd206, 8'd41, 1'b1, 1'b0};
2070: data_out = {8'd207, 8'd41, 1'b1, 1'b0};
2071: data_out = {8'd208, 8'd41, 1'b1, 1'b0};
2072: data_out = {8'd209, 8'd41, 1'b1, 1'b0};
2073: data_out = {8'd210, 8'd41, 1'b1, 1'b0};
2074: data_out = {8'd211, 8'd41, 1'b1, 1'b0};
2075: data_out = {8'd6, 8'd42, 1'b1, 1'b0};
2076: data_out = {8'd7, 8'd42, 1'b1, 1'b0};
2077: data_out = {8'd8, 8'd42, 1'b1, 1'b0};
2078: data_out = {8'd9, 8'd42, 1'b1, 1'b0};
2079: data_out = {8'd10, 8'd42, 1'b1, 1'b0};
2080: data_out = {8'd11, 8'd42, 1'b1, 1'b0};
2081: data_out = {8'd25, 8'd42, 1'b1, 1'b0};
2082: data_out = {8'd26, 8'd42, 1'b1, 1'b0};
2083: data_out = {8'd27, 8'd42, 1'b1, 1'b0};
2084: data_out = {8'd28, 8'd42, 1'b1, 1'b0};
2085: data_out = {8'd29, 8'd42, 1'b1, 1'b0};
2086: data_out = {8'd30, 8'd42, 1'b1, 1'b0};
2087: data_out = {8'd36, 8'd42, 1'b1, 1'b0};
2088: data_out = {8'd37, 8'd42, 1'b1, 1'b0};
2089: data_out = {8'd38, 8'd42, 1'b1, 1'b0};
2090: data_out = {8'd39, 8'd42, 1'b1, 1'b0};
2091: data_out = {8'd40, 8'd42, 1'b1, 1'b0};
2092: data_out = {8'd41, 8'd42, 1'b1, 1'b0};
2093: data_out = {8'd55, 8'd42, 1'b1, 1'b0};
2094: data_out = {8'd56, 8'd42, 1'b1, 1'b0};
2095: data_out = {8'd57, 8'd42, 1'b1, 1'b0};
2096: data_out = {8'd58, 8'd42, 1'b1, 1'b0};
2097: data_out = {8'd59, 8'd42, 1'b1, 1'b0};
2098: data_out = {8'd60, 8'd42, 1'b1, 1'b0};
2099: data_out = {8'd73, 8'd42, 1'b1, 1'b0};
2100: data_out = {8'd74, 8'd42, 1'b1, 1'b0};
2101: data_out = {8'd75, 8'd42, 1'b1, 1'b0};
2102: data_out = {8'd76, 8'd42, 1'b1, 1'b0};
2103: data_out = {8'd77, 8'd42, 1'b1, 1'b0};
2104: data_out = {8'd78, 8'd42, 1'b1, 1'b0};
2105: data_out = {8'd97, 8'd42, 1'b1, 1'b0};
2106: data_out = {8'd98, 8'd42, 1'b1, 1'b0};
2107: data_out = {8'd99, 8'd42, 1'b1, 1'b0};
2108: data_out = {8'd100, 8'd42, 1'b1, 1'b0};
2109: data_out = {8'd101, 8'd42, 1'b1, 1'b0};
2110: data_out = {8'd102, 8'd42, 1'b1, 1'b0};
2111: data_out = {8'd116, 8'd42, 1'b1, 1'b0};
2112: data_out = {8'd117, 8'd42, 1'b1, 1'b0};
2113: data_out = {8'd118, 8'd42, 1'b1, 1'b0};
2114: data_out = {8'd119, 8'd42, 1'b1, 1'b0};
2115: data_out = {8'd120, 8'd42, 1'b1, 1'b0};
2116: data_out = {8'd121, 8'd42, 1'b1, 1'b0};
2117: data_out = {8'd127, 8'd42, 1'b1, 1'b0};
2118: data_out = {8'd128, 8'd42, 1'b1, 1'b0};
2119: data_out = {8'd129, 8'd42, 1'b1, 1'b0};
2120: data_out = {8'd130, 8'd42, 1'b1, 1'b0};
2121: data_out = {8'd131, 8'd42, 1'b1, 1'b0};
2122: data_out = {8'd132, 8'd42, 1'b1, 1'b0};
2123: data_out = {8'd146, 8'd42, 1'b1, 1'b0};
2124: data_out = {8'd147, 8'd42, 1'b1, 1'b0};
2125: data_out = {8'd148, 8'd42, 1'b1, 1'b0};
2126: data_out = {8'd149, 8'd42, 1'b1, 1'b0};
2127: data_out = {8'd150, 8'd42, 1'b1, 1'b0};
2128: data_out = {8'd151, 8'd42, 1'b1, 1'b0};
2129: data_out = {8'd187, 8'd42, 1'b1, 1'b0};
2130: data_out = {8'd188, 8'd42, 1'b1, 1'b0};
2131: data_out = {8'd189, 8'd42, 1'b1, 1'b0};
2132: data_out = {8'd190, 8'd42, 1'b1, 1'b0};
2133: data_out = {8'd191, 8'd42, 1'b1, 1'b0};
2134: data_out = {8'd192, 8'd42, 1'b1, 1'b0};
2135: data_out = {8'd206, 8'd42, 1'b1, 1'b0};
2136: data_out = {8'd207, 8'd42, 1'b1, 1'b0};
2137: data_out = {8'd208, 8'd42, 1'b1, 1'b0};
2138: data_out = {8'd209, 8'd42, 1'b1, 1'b0};
2139: data_out = {8'd210, 8'd42, 1'b1, 1'b0};
2140: data_out = {8'd211, 8'd42, 1'b1, 1'b0};
2141: data_out = {8'd6, 8'd43, 1'b1, 1'b0};
2142: data_out = {8'd7, 8'd43, 1'b1, 1'b0};
2143: data_out = {8'd8, 8'd43, 1'b1, 1'b0};
2144: data_out = {8'd9, 8'd43, 1'b1, 1'b0};
2145: data_out = {8'd10, 8'd43, 1'b1, 1'b0};
2146: data_out = {8'd11, 8'd43, 1'b1, 1'b0};
2147: data_out = {8'd25, 8'd43, 1'b1, 1'b0};
2148: data_out = {8'd26, 8'd43, 1'b1, 1'b0};
2149: data_out = {8'd27, 8'd43, 1'b1, 1'b0};
2150: data_out = {8'd28, 8'd43, 1'b1, 1'b0};
2151: data_out = {8'd29, 8'd43, 1'b1, 1'b0};
2152: data_out = {8'd30, 8'd43, 1'b1, 1'b0};
2153: data_out = {8'd36, 8'd43, 1'b1, 1'b0};
2154: data_out = {8'd37, 8'd43, 1'b1, 1'b0};
2155: data_out = {8'd38, 8'd43, 1'b1, 1'b0};
2156: data_out = {8'd39, 8'd43, 1'b1, 1'b0};
2157: data_out = {8'd40, 8'd43, 1'b1, 1'b0};
2158: data_out = {8'd41, 8'd43, 1'b1, 1'b0};
2159: data_out = {8'd55, 8'd43, 1'b1, 1'b0};
2160: data_out = {8'd56, 8'd43, 1'b1, 1'b0};
2161: data_out = {8'd57, 8'd43, 1'b1, 1'b0};
2162: data_out = {8'd58, 8'd43, 1'b1, 1'b0};
2163: data_out = {8'd59, 8'd43, 1'b1, 1'b0};
2164: data_out = {8'd60, 8'd43, 1'b1, 1'b0};
2165: data_out = {8'd73, 8'd43, 1'b1, 1'b0};
2166: data_out = {8'd74, 8'd43, 1'b1, 1'b0};
2167: data_out = {8'd75, 8'd43, 1'b1, 1'b0};
2168: data_out = {8'd76, 8'd43, 1'b1, 1'b0};
2169: data_out = {8'd77, 8'd43, 1'b1, 1'b0};
2170: data_out = {8'd78, 8'd43, 1'b1, 1'b0};
2171: data_out = {8'd97, 8'd43, 1'b1, 1'b0};
2172: data_out = {8'd98, 8'd43, 1'b1, 1'b0};
2173: data_out = {8'd99, 8'd43, 1'b1, 1'b0};
2174: data_out = {8'd100, 8'd43, 1'b1, 1'b0};
2175: data_out = {8'd101, 8'd43, 1'b1, 1'b0};
2176: data_out = {8'd102, 8'd43, 1'b1, 1'b0};
2177: data_out = {8'd116, 8'd43, 1'b1, 1'b0};
2178: data_out = {8'd117, 8'd43, 1'b1, 1'b0};
2179: data_out = {8'd118, 8'd43, 1'b1, 1'b0};
2180: data_out = {8'd119, 8'd43, 1'b1, 1'b0};
2181: data_out = {8'd120, 8'd43, 1'b1, 1'b0};
2182: data_out = {8'd121, 8'd43, 1'b1, 1'b0};
2183: data_out = {8'd127, 8'd43, 1'b1, 1'b0};
2184: data_out = {8'd128, 8'd43, 1'b1, 1'b0};
2185: data_out = {8'd129, 8'd43, 1'b1, 1'b0};
2186: data_out = {8'd130, 8'd43, 1'b1, 1'b0};
2187: data_out = {8'd131, 8'd43, 1'b1, 1'b0};
2188: data_out = {8'd132, 8'd43, 1'b1, 1'b0};
2189: data_out = {8'd146, 8'd43, 1'b1, 1'b0};
2190: data_out = {8'd147, 8'd43, 1'b1, 1'b0};
2191: data_out = {8'd148, 8'd43, 1'b1, 1'b0};
2192: data_out = {8'd149, 8'd43, 1'b1, 1'b0};
2193: data_out = {8'd150, 8'd43, 1'b1, 1'b0};
2194: data_out = {8'd151, 8'd43, 1'b1, 1'b0};
2195: data_out = {8'd187, 8'd43, 1'b1, 1'b0};
2196: data_out = {8'd188, 8'd43, 1'b1, 1'b0};
2197: data_out = {8'd189, 8'd43, 1'b1, 1'b0};
2198: data_out = {8'd190, 8'd43, 1'b1, 1'b0};
2199: data_out = {8'd191, 8'd43, 1'b1, 1'b0};
2200: data_out = {8'd192, 8'd43, 1'b1, 1'b0};
2201: data_out = {8'd206, 8'd43, 1'b1, 1'b0};
2202: data_out = {8'd207, 8'd43, 1'b1, 1'b0};
2203: data_out = {8'd208, 8'd43, 1'b1, 1'b0};
2204: data_out = {8'd209, 8'd43, 1'b1, 1'b0};
2205: data_out = {8'd210, 8'd43, 1'b1, 1'b0};
2206: data_out = {8'd211, 8'd43, 1'b1, 1'b0};
2207: data_out = {8'd6, 8'd44, 1'b1, 1'b0};
2208: data_out = {8'd7, 8'd44, 1'b1, 1'b0};
2209: data_out = {8'd8, 8'd44, 1'b1, 1'b0};
2210: data_out = {8'd9, 8'd44, 1'b1, 1'b0};
2211: data_out = {8'd10, 8'd44, 1'b1, 1'b0};
2212: data_out = {8'd11, 8'd44, 1'b1, 1'b0};
2213: data_out = {8'd25, 8'd44, 1'b1, 1'b0};
2214: data_out = {8'd26, 8'd44, 1'b1, 1'b0};
2215: data_out = {8'd27, 8'd44, 1'b1, 1'b0};
2216: data_out = {8'd28, 8'd44, 1'b1, 1'b0};
2217: data_out = {8'd29, 8'd44, 1'b1, 1'b0};
2218: data_out = {8'd30, 8'd44, 1'b1, 1'b0};
2219: data_out = {8'd36, 8'd44, 1'b1, 1'b0};
2220: data_out = {8'd37, 8'd44, 1'b1, 1'b0};
2221: data_out = {8'd38, 8'd44, 1'b1, 1'b0};
2222: data_out = {8'd39, 8'd44, 1'b1, 1'b0};
2223: data_out = {8'd40, 8'd44, 1'b1, 1'b0};
2224: data_out = {8'd41, 8'd44, 1'b1, 1'b0};
2225: data_out = {8'd55, 8'd44, 1'b1, 1'b0};
2226: data_out = {8'd56, 8'd44, 1'b1, 1'b0};
2227: data_out = {8'd57, 8'd44, 1'b1, 1'b0};
2228: data_out = {8'd58, 8'd44, 1'b1, 1'b0};
2229: data_out = {8'd59, 8'd44, 1'b1, 1'b0};
2230: data_out = {8'd60, 8'd44, 1'b1, 1'b0};
2231: data_out = {8'd73, 8'd44, 1'b1, 1'b0};
2232: data_out = {8'd74, 8'd44, 1'b1, 1'b0};
2233: data_out = {8'd75, 8'd44, 1'b1, 1'b0};
2234: data_out = {8'd76, 8'd44, 1'b1, 1'b0};
2235: data_out = {8'd77, 8'd44, 1'b1, 1'b0};
2236: data_out = {8'd78, 8'd44, 1'b1, 1'b0};
2237: data_out = {8'd97, 8'd44, 1'b1, 1'b0};
2238: data_out = {8'd98, 8'd44, 1'b1, 1'b0};
2239: data_out = {8'd99, 8'd44, 1'b1, 1'b0};
2240: data_out = {8'd100, 8'd44, 1'b1, 1'b0};
2241: data_out = {8'd101, 8'd44, 1'b1, 1'b0};
2242: data_out = {8'd102, 8'd44, 1'b1, 1'b0};
2243: data_out = {8'd116, 8'd44, 1'b1, 1'b0};
2244: data_out = {8'd117, 8'd44, 1'b1, 1'b0};
2245: data_out = {8'd118, 8'd44, 1'b1, 1'b0};
2246: data_out = {8'd119, 8'd44, 1'b1, 1'b0};
2247: data_out = {8'd120, 8'd44, 1'b1, 1'b0};
2248: data_out = {8'd121, 8'd44, 1'b1, 1'b0};
2249: data_out = {8'd127, 8'd44, 1'b1, 1'b0};
2250: data_out = {8'd128, 8'd44, 1'b1, 1'b0};
2251: data_out = {8'd129, 8'd44, 1'b1, 1'b0};
2252: data_out = {8'd130, 8'd44, 1'b1, 1'b0};
2253: data_out = {8'd131, 8'd44, 1'b1, 1'b0};
2254: data_out = {8'd132, 8'd44, 1'b1, 1'b0};
2255: data_out = {8'd146, 8'd44, 1'b1, 1'b0};
2256: data_out = {8'd147, 8'd44, 1'b1, 1'b0};
2257: data_out = {8'd148, 8'd44, 1'b1, 1'b0};
2258: data_out = {8'd149, 8'd44, 1'b1, 1'b0};
2259: data_out = {8'd150, 8'd44, 1'b1, 1'b0};
2260: data_out = {8'd151, 8'd44, 1'b1, 1'b0};
2261: data_out = {8'd187, 8'd44, 1'b1, 1'b0};
2262: data_out = {8'd188, 8'd44, 1'b1, 1'b0};
2263: data_out = {8'd189, 8'd44, 1'b1, 1'b0};
2264: data_out = {8'd190, 8'd44, 1'b1, 1'b0};
2265: data_out = {8'd191, 8'd44, 1'b1, 1'b0};
2266: data_out = {8'd192, 8'd44, 1'b1, 1'b0};
2267: data_out = {8'd206, 8'd44, 1'b1, 1'b0};
2268: data_out = {8'd207, 8'd44, 1'b1, 1'b0};
2269: data_out = {8'd208, 8'd44, 1'b1, 1'b0};
2270: data_out = {8'd209, 8'd44, 1'b1, 1'b0};
2271: data_out = {8'd210, 8'd44, 1'b1, 1'b0};
2272: data_out = {8'd211, 8'd44, 1'b1, 1'b0};
2273: data_out = {8'd6, 8'd45, 1'b1, 1'b0};
2274: data_out = {8'd7, 8'd45, 1'b1, 1'b0};
2275: data_out = {8'd8, 8'd45, 1'b1, 1'b0};
2276: data_out = {8'd9, 8'd45, 1'b1, 1'b0};
2277: data_out = {8'd10, 8'd45, 1'b1, 1'b0};
2278: data_out = {8'd11, 8'd45, 1'b1, 1'b0};
2279: data_out = {8'd25, 8'd45, 1'b1, 1'b0};
2280: data_out = {8'd26, 8'd45, 1'b1, 1'b0};
2281: data_out = {8'd27, 8'd45, 1'b1, 1'b0};
2282: data_out = {8'd28, 8'd45, 1'b1, 1'b0};
2283: data_out = {8'd29, 8'd45, 1'b1, 1'b0};
2284: data_out = {8'd30, 8'd45, 1'b1, 1'b0};
2285: data_out = {8'd36, 8'd45, 1'b1, 1'b0};
2286: data_out = {8'd37, 8'd45, 1'b1, 1'b0};
2287: data_out = {8'd38, 8'd45, 1'b1, 1'b0};
2288: data_out = {8'd39, 8'd45, 1'b1, 1'b0};
2289: data_out = {8'd40, 8'd45, 1'b1, 1'b0};
2290: data_out = {8'd41, 8'd45, 1'b1, 1'b0};
2291: data_out = {8'd55, 8'd45, 1'b1, 1'b0};
2292: data_out = {8'd56, 8'd45, 1'b1, 1'b0};
2293: data_out = {8'd57, 8'd45, 1'b1, 1'b0};
2294: data_out = {8'd58, 8'd45, 1'b1, 1'b0};
2295: data_out = {8'd59, 8'd45, 1'b1, 1'b0};
2296: data_out = {8'd60, 8'd45, 1'b1, 1'b0};
2297: data_out = {8'd73, 8'd45, 1'b1, 1'b0};
2298: data_out = {8'd74, 8'd45, 1'b1, 1'b0};
2299: data_out = {8'd75, 8'd45, 1'b1, 1'b0};
2300: data_out = {8'd76, 8'd45, 1'b1, 1'b0};
2301: data_out = {8'd77, 8'd45, 1'b1, 1'b0};
2302: data_out = {8'd78, 8'd45, 1'b1, 1'b0};
2303: data_out = {8'd97, 8'd45, 1'b1, 1'b0};
2304: data_out = {8'd98, 8'd45, 1'b1, 1'b0};
2305: data_out = {8'd99, 8'd45, 1'b1, 1'b0};
2306: data_out = {8'd100, 8'd45, 1'b1, 1'b0};
2307: data_out = {8'd101, 8'd45, 1'b1, 1'b0};
2308: data_out = {8'd102, 8'd45, 1'b1, 1'b0};
2309: data_out = {8'd116, 8'd45, 1'b1, 1'b0};
2310: data_out = {8'd117, 8'd45, 1'b1, 1'b0};
2311: data_out = {8'd118, 8'd45, 1'b1, 1'b0};
2312: data_out = {8'd119, 8'd45, 1'b1, 1'b0};
2313: data_out = {8'd120, 8'd45, 1'b1, 1'b0};
2314: data_out = {8'd121, 8'd45, 1'b1, 1'b0};
2315: data_out = {8'd127, 8'd45, 1'b1, 1'b0};
2316: data_out = {8'd128, 8'd45, 1'b1, 1'b0};
2317: data_out = {8'd129, 8'd45, 1'b1, 1'b0};
2318: data_out = {8'd130, 8'd45, 1'b1, 1'b0};
2319: data_out = {8'd131, 8'd45, 1'b1, 1'b0};
2320: data_out = {8'd132, 8'd45, 1'b1, 1'b0};
2321: data_out = {8'd146, 8'd45, 1'b1, 1'b0};
2322: data_out = {8'd147, 8'd45, 1'b1, 1'b0};
2323: data_out = {8'd148, 8'd45, 1'b1, 1'b0};
2324: data_out = {8'd149, 8'd45, 1'b1, 1'b0};
2325: data_out = {8'd150, 8'd45, 1'b1, 1'b0};
2326: data_out = {8'd151, 8'd45, 1'b1, 1'b0};
2327: data_out = {8'd187, 8'd45, 1'b1, 1'b0};
2328: data_out = {8'd188, 8'd45, 1'b1, 1'b0};
2329: data_out = {8'd189, 8'd45, 1'b1, 1'b0};
2330: data_out = {8'd190, 8'd45, 1'b1, 1'b0};
2331: data_out = {8'd191, 8'd45, 1'b1, 1'b0};
2332: data_out = {8'd192, 8'd45, 1'b1, 1'b0};
2333: data_out = {8'd206, 8'd45, 1'b1, 1'b0};
2334: data_out = {8'd207, 8'd45, 1'b1, 1'b0};
2335: data_out = {8'd208, 8'd45, 1'b1, 1'b0};
2336: data_out = {8'd209, 8'd45, 1'b1, 1'b0};
2337: data_out = {8'd210, 8'd45, 1'b1, 1'b0};
2338: data_out = {8'd211, 8'd45, 1'b1, 1'b0};
2339: data_out = {8'd6, 8'd46, 1'b1, 1'b0};
2340: data_out = {8'd7, 8'd46, 1'b1, 1'b0};
2341: data_out = {8'd8, 8'd46, 1'b1, 1'b0};
2342: data_out = {8'd9, 8'd46, 1'b1, 1'b0};
2343: data_out = {8'd10, 8'd46, 1'b1, 1'b0};
2344: data_out = {8'd11, 8'd46, 1'b1, 1'b0};
2345: data_out = {8'd25, 8'd46, 1'b1, 1'b0};
2346: data_out = {8'd26, 8'd46, 1'b1, 1'b0};
2347: data_out = {8'd27, 8'd46, 1'b1, 1'b0};
2348: data_out = {8'd28, 8'd46, 1'b1, 1'b0};
2349: data_out = {8'd29, 8'd46, 1'b1, 1'b0};
2350: data_out = {8'd30, 8'd46, 1'b1, 1'b0};
2351: data_out = {8'd36, 8'd46, 1'b1, 1'b0};
2352: data_out = {8'd37, 8'd46, 1'b1, 1'b0};
2353: data_out = {8'd38, 8'd46, 1'b1, 1'b0};
2354: data_out = {8'd39, 8'd46, 1'b1, 1'b0};
2355: data_out = {8'd40, 8'd46, 1'b1, 1'b0};
2356: data_out = {8'd41, 8'd46, 1'b1, 1'b0};
2357: data_out = {8'd55, 8'd46, 1'b1, 1'b0};
2358: data_out = {8'd56, 8'd46, 1'b1, 1'b0};
2359: data_out = {8'd57, 8'd46, 1'b1, 1'b0};
2360: data_out = {8'd58, 8'd46, 1'b1, 1'b0};
2361: data_out = {8'd59, 8'd46, 1'b1, 1'b0};
2362: data_out = {8'd60, 8'd46, 1'b1, 1'b0};
2363: data_out = {8'd73, 8'd46, 1'b1, 1'b0};
2364: data_out = {8'd74, 8'd46, 1'b1, 1'b0};
2365: data_out = {8'd75, 8'd46, 1'b1, 1'b0};
2366: data_out = {8'd76, 8'd46, 1'b1, 1'b0};
2367: data_out = {8'd77, 8'd46, 1'b1, 1'b0};
2368: data_out = {8'd78, 8'd46, 1'b1, 1'b0};
2369: data_out = {8'd97, 8'd46, 1'b1, 1'b0};
2370: data_out = {8'd98, 8'd46, 1'b1, 1'b0};
2371: data_out = {8'd99, 8'd46, 1'b1, 1'b0};
2372: data_out = {8'd100, 8'd46, 1'b1, 1'b0};
2373: data_out = {8'd101, 8'd46, 1'b1, 1'b0};
2374: data_out = {8'd102, 8'd46, 1'b1, 1'b0};
2375: data_out = {8'd116, 8'd46, 1'b1, 1'b0};
2376: data_out = {8'd117, 8'd46, 1'b1, 1'b0};
2377: data_out = {8'd118, 8'd46, 1'b1, 1'b0};
2378: data_out = {8'd119, 8'd46, 1'b1, 1'b0};
2379: data_out = {8'd120, 8'd46, 1'b1, 1'b0};
2380: data_out = {8'd121, 8'd46, 1'b1, 1'b0};
2381: data_out = {8'd127, 8'd46, 1'b1, 1'b0};
2382: data_out = {8'd128, 8'd46, 1'b1, 1'b0};
2383: data_out = {8'd129, 8'd46, 1'b1, 1'b0};
2384: data_out = {8'd130, 8'd46, 1'b1, 1'b0};
2385: data_out = {8'd131, 8'd46, 1'b1, 1'b0};
2386: data_out = {8'd132, 8'd46, 1'b1, 1'b0};
2387: data_out = {8'd146, 8'd46, 1'b1, 1'b0};
2388: data_out = {8'd147, 8'd46, 1'b1, 1'b0};
2389: data_out = {8'd148, 8'd46, 1'b1, 1'b0};
2390: data_out = {8'd149, 8'd46, 1'b1, 1'b0};
2391: data_out = {8'd150, 8'd46, 1'b1, 1'b0};
2392: data_out = {8'd151, 8'd46, 1'b1, 1'b0};
2393: data_out = {8'd187, 8'd46, 1'b1, 1'b0};
2394: data_out = {8'd188, 8'd46, 1'b1, 1'b0};
2395: data_out = {8'd189, 8'd46, 1'b1, 1'b0};
2396: data_out = {8'd190, 8'd46, 1'b1, 1'b0};
2397: data_out = {8'd191, 8'd46, 1'b1, 1'b0};
2398: data_out = {8'd192, 8'd46, 1'b1, 1'b0};
2399: data_out = {8'd206, 8'd46, 1'b1, 1'b0};
2400: data_out = {8'd207, 8'd46, 1'b1, 1'b0};
2401: data_out = {8'd208, 8'd46, 1'b1, 1'b0};
2402: data_out = {8'd209, 8'd46, 1'b1, 1'b0};
2403: data_out = {8'd210, 8'd46, 1'b1, 1'b0};
2404: data_out = {8'd211, 8'd46, 1'b1, 1'b0};
2405: data_out = {8'd6, 8'd47, 1'b1, 1'b0};
2406: data_out = {8'd7, 8'd47, 1'b1, 1'b0};
2407: data_out = {8'd8, 8'd47, 1'b1, 1'b0};
2408: data_out = {8'd9, 8'd47, 1'b1, 1'b0};
2409: data_out = {8'd10, 8'd47, 1'b1, 1'b0};
2410: data_out = {8'd11, 8'd47, 1'b1, 1'b0};
2411: data_out = {8'd25, 8'd47, 1'b1, 1'b0};
2412: data_out = {8'd26, 8'd47, 1'b1, 1'b0};
2413: data_out = {8'd27, 8'd47, 1'b1, 1'b0};
2414: data_out = {8'd28, 8'd47, 1'b1, 1'b0};
2415: data_out = {8'd29, 8'd47, 1'b1, 1'b0};
2416: data_out = {8'd30, 8'd47, 1'b1, 1'b0};
2417: data_out = {8'd36, 8'd47, 1'b1, 1'b0};
2418: data_out = {8'd37, 8'd47, 1'b1, 1'b0};
2419: data_out = {8'd38, 8'd47, 1'b1, 1'b0};
2420: data_out = {8'd39, 8'd47, 1'b1, 1'b0};
2421: data_out = {8'd40, 8'd47, 1'b1, 1'b0};
2422: data_out = {8'd41, 8'd47, 1'b1, 1'b0};
2423: data_out = {8'd55, 8'd47, 1'b1, 1'b0};
2424: data_out = {8'd56, 8'd47, 1'b1, 1'b0};
2425: data_out = {8'd57, 8'd47, 1'b1, 1'b0};
2426: data_out = {8'd58, 8'd47, 1'b1, 1'b0};
2427: data_out = {8'd59, 8'd47, 1'b1, 1'b0};
2428: data_out = {8'd60, 8'd47, 1'b1, 1'b0};
2429: data_out = {8'd73, 8'd47, 1'b1, 1'b0};
2430: data_out = {8'd74, 8'd47, 1'b1, 1'b0};
2431: data_out = {8'd75, 8'd47, 1'b1, 1'b0};
2432: data_out = {8'd76, 8'd47, 1'b1, 1'b0};
2433: data_out = {8'd77, 8'd47, 1'b1, 1'b0};
2434: data_out = {8'd78, 8'd47, 1'b1, 1'b0};
2435: data_out = {8'd97, 8'd47, 1'b1, 1'b0};
2436: data_out = {8'd98, 8'd47, 1'b1, 1'b0};
2437: data_out = {8'd99, 8'd47, 1'b1, 1'b0};
2438: data_out = {8'd100, 8'd47, 1'b1, 1'b0};
2439: data_out = {8'd101, 8'd47, 1'b1, 1'b0};
2440: data_out = {8'd102, 8'd47, 1'b1, 1'b0};
2441: data_out = {8'd116, 8'd47, 1'b1, 1'b0};
2442: data_out = {8'd117, 8'd47, 1'b1, 1'b0};
2443: data_out = {8'd118, 8'd47, 1'b1, 1'b0};
2444: data_out = {8'd119, 8'd47, 1'b1, 1'b0};
2445: data_out = {8'd120, 8'd47, 1'b1, 1'b0};
2446: data_out = {8'd121, 8'd47, 1'b1, 1'b0};
2447: data_out = {8'd127, 8'd47, 1'b1, 1'b0};
2448: data_out = {8'd128, 8'd47, 1'b1, 1'b0};
2449: data_out = {8'd129, 8'd47, 1'b1, 1'b0};
2450: data_out = {8'd130, 8'd47, 1'b1, 1'b0};
2451: data_out = {8'd131, 8'd47, 1'b1, 1'b0};
2452: data_out = {8'd132, 8'd47, 1'b1, 1'b0};
2453: data_out = {8'd146, 8'd47, 1'b1, 1'b0};
2454: data_out = {8'd147, 8'd47, 1'b1, 1'b0};
2455: data_out = {8'd148, 8'd47, 1'b1, 1'b0};
2456: data_out = {8'd149, 8'd47, 1'b1, 1'b0};
2457: data_out = {8'd150, 8'd47, 1'b1, 1'b0};
2458: data_out = {8'd151, 8'd47, 1'b1, 1'b0};
2459: data_out = {8'd187, 8'd47, 1'b1, 1'b0};
2460: data_out = {8'd188, 8'd47, 1'b1, 1'b0};
2461: data_out = {8'd189, 8'd47, 1'b1, 1'b0};
2462: data_out = {8'd190, 8'd47, 1'b1, 1'b0};
2463: data_out = {8'd191, 8'd47, 1'b1, 1'b0};
2464: data_out = {8'd192, 8'd47, 1'b1, 1'b0};
2465: data_out = {8'd206, 8'd47, 1'b1, 1'b0};
2466: data_out = {8'd207, 8'd47, 1'b1, 1'b0};
2467: data_out = {8'd208, 8'd47, 1'b1, 1'b0};
2468: data_out = {8'd209, 8'd47, 1'b1, 1'b0};
2469: data_out = {8'd210, 8'd47, 1'b1, 1'b0};
2470: data_out = {8'd211, 8'd47, 1'b1, 1'b0};
2471: data_out = {8'd6, 8'd48, 1'b1, 1'b0};
2472: data_out = {8'd7, 8'd48, 1'b1, 1'b0};
2473: data_out = {8'd8, 8'd48, 1'b1, 1'b0};
2474: data_out = {8'd9, 8'd48, 1'b1, 1'b0};
2475: data_out = {8'd10, 8'd48, 1'b1, 1'b0};
2476: data_out = {8'd11, 8'd48, 1'b1, 1'b0};
2477: data_out = {8'd25, 8'd48, 1'b1, 1'b0};
2478: data_out = {8'd26, 8'd48, 1'b1, 1'b0};
2479: data_out = {8'd27, 8'd48, 1'b1, 1'b0};
2480: data_out = {8'd28, 8'd48, 1'b1, 1'b0};
2481: data_out = {8'd29, 8'd48, 1'b1, 1'b0};
2482: data_out = {8'd30, 8'd48, 1'b1, 1'b0};
2483: data_out = {8'd36, 8'd48, 1'b1, 1'b0};
2484: data_out = {8'd37, 8'd48, 1'b1, 1'b0};
2485: data_out = {8'd38, 8'd48, 1'b1, 1'b0};
2486: data_out = {8'd39, 8'd48, 1'b1, 1'b0};
2487: data_out = {8'd40, 8'd48, 1'b1, 1'b0};
2488: data_out = {8'd41, 8'd48, 1'b1, 1'b0};
2489: data_out = {8'd42, 8'd48, 1'b1, 1'b0};
2490: data_out = {8'd43, 8'd48, 1'b1, 1'b0};
2491: data_out = {8'd44, 8'd48, 1'b1, 1'b0};
2492: data_out = {8'd45, 8'd48, 1'b1, 1'b0};
2493: data_out = {8'd46, 8'd48, 1'b1, 1'b0};
2494: data_out = {8'd47, 8'd48, 1'b1, 1'b0};
2495: data_out = {8'd48, 8'd48, 1'b1, 1'b0};
2496: data_out = {8'd49, 8'd48, 1'b1, 1'b0};
2497: data_out = {8'd50, 8'd48, 1'b1, 1'b0};
2498: data_out = {8'd51, 8'd48, 1'b1, 1'b0};
2499: data_out = {8'd52, 8'd48, 1'b1, 1'b0};
2500: data_out = {8'd53, 8'd48, 1'b1, 1'b0};
2501: data_out = {8'd54, 8'd48, 1'b1, 1'b0};
2502: data_out = {8'd55, 8'd48, 1'b1, 1'b0};
2503: data_out = {8'd56, 8'd48, 1'b1, 1'b0};
2504: data_out = {8'd57, 8'd48, 1'b1, 1'b0};
2505: data_out = {8'd58, 8'd48, 1'b1, 1'b0};
2506: data_out = {8'd59, 8'd48, 1'b1, 1'b0};
2507: data_out = {8'd60, 8'd48, 1'b1, 1'b0};
2508: data_out = {8'd63, 8'd48, 1'b1, 1'b0};
2509: data_out = {8'd64, 8'd48, 1'b1, 1'b0};
2510: data_out = {8'd65, 8'd48, 1'b1, 1'b0};
2511: data_out = {8'd66, 8'd48, 1'b1, 1'b0};
2512: data_out = {8'd67, 8'd48, 1'b1, 1'b0};
2513: data_out = {8'd68, 8'd48, 1'b1, 1'b0};
2514: data_out = {8'd69, 8'd48, 1'b1, 1'b0};
2515: data_out = {8'd70, 8'd48, 1'b1, 1'b0};
2516: data_out = {8'd71, 8'd48, 1'b1, 1'b0};
2517: data_out = {8'd72, 8'd48, 1'b1, 1'b0};
2518: data_out = {8'd73, 8'd48, 1'b1, 1'b0};
2519: data_out = {8'd74, 8'd48, 1'b1, 1'b0};
2520: data_out = {8'd75, 8'd48, 1'b1, 1'b0};
2521: data_out = {8'd76, 8'd48, 1'b1, 1'b0};
2522: data_out = {8'd77, 8'd48, 1'b1, 1'b0};
2523: data_out = {8'd78, 8'd48, 1'b1, 1'b0};
2524: data_out = {8'd79, 8'd48, 1'b1, 1'b0};
2525: data_out = {8'd80, 8'd48, 1'b1, 1'b0};
2526: data_out = {8'd81, 8'd48, 1'b1, 1'b0};
2527: data_out = {8'd82, 8'd48, 1'b1, 1'b0};
2528: data_out = {8'd83, 8'd48, 1'b1, 1'b0};
2529: data_out = {8'd84, 8'd48, 1'b1, 1'b0};
2530: data_out = {8'd85, 8'd48, 1'b1, 1'b0};
2531: data_out = {8'd86, 8'd48, 1'b1, 1'b0};
2532: data_out = {8'd87, 8'd48, 1'b1, 1'b0};
2533: data_out = {8'd88, 8'd48, 1'b1, 1'b0};
2534: data_out = {8'd89, 8'd48, 1'b1, 1'b0};
2535: data_out = {8'd90, 8'd48, 1'b1, 1'b0};
2536: data_out = {8'd91, 8'd48, 1'b1, 1'b0};
2537: data_out = {8'd97, 8'd48, 1'b1, 1'b0};
2538: data_out = {8'd98, 8'd48, 1'b1, 1'b0};
2539: data_out = {8'd99, 8'd48, 1'b1, 1'b0};
2540: data_out = {8'd100, 8'd48, 1'b1, 1'b0};
2541: data_out = {8'd101, 8'd48, 1'b1, 1'b0};
2542: data_out = {8'd102, 8'd48, 1'b1, 1'b0};
2543: data_out = {8'd103, 8'd48, 1'b1, 1'b0};
2544: data_out = {8'd104, 8'd48, 1'b1, 1'b0};
2545: data_out = {8'd105, 8'd48, 1'b1, 1'b0};
2546: data_out = {8'd106, 8'd48, 1'b1, 1'b0};
2547: data_out = {8'd107, 8'd48, 1'b1, 1'b0};
2548: data_out = {8'd108, 8'd48, 1'b1, 1'b0};
2549: data_out = {8'd109, 8'd48, 1'b1, 1'b0};
2550: data_out = {8'd110, 8'd48, 1'b1, 1'b0};
2551: data_out = {8'd111, 8'd48, 1'b1, 1'b0};
2552: data_out = {8'd112, 8'd48, 1'b1, 1'b0};
2553: data_out = {8'd113, 8'd48, 1'b1, 1'b0};
2554: data_out = {8'd114, 8'd48, 1'b1, 1'b0};
2555: data_out = {8'd115, 8'd48, 1'b1, 1'b0};
2556: data_out = {8'd116, 8'd48, 1'b1, 1'b0};
2557: data_out = {8'd117, 8'd48, 1'b1, 1'b0};
2558: data_out = {8'd118, 8'd48, 1'b1, 1'b0};
2559: data_out = {8'd119, 8'd48, 1'b1, 1'b0};
2560: data_out = {8'd120, 8'd48, 1'b1, 1'b0};
2561: data_out = {8'd121, 8'd48, 1'b1, 1'b0};
2562: data_out = {8'd127, 8'd48, 1'b1, 1'b0};
2563: data_out = {8'd128, 8'd48, 1'b1, 1'b0};
2564: data_out = {8'd129, 8'd48, 1'b1, 1'b0};
2565: data_out = {8'd130, 8'd48, 1'b1, 1'b0};
2566: data_out = {8'd131, 8'd48, 1'b1, 1'b0};
2567: data_out = {8'd132, 8'd48, 1'b1, 1'b0};
2568: data_out = {8'd133, 8'd48, 1'b1, 1'b0};
2569: data_out = {8'd134, 8'd48, 1'b1, 1'b0};
2570: data_out = {8'd135, 8'd48, 1'b1, 1'b0};
2571: data_out = {8'd136, 8'd48, 1'b1, 1'b0};
2572: data_out = {8'd137, 8'd48, 1'b1, 1'b0};
2573: data_out = {8'd138, 8'd48, 1'b1, 1'b0};
2574: data_out = {8'd139, 8'd48, 1'b1, 1'b0};
2575: data_out = {8'd140, 8'd48, 1'b1, 1'b0};
2576: data_out = {8'd141, 8'd48, 1'b1, 1'b0};
2577: data_out = {8'd142, 8'd48, 1'b1, 1'b0};
2578: data_out = {8'd143, 8'd48, 1'b1, 1'b0};
2579: data_out = {8'd144, 8'd48, 1'b1, 1'b0};
2580: data_out = {8'd145, 8'd48, 1'b1, 1'b0};
2581: data_out = {8'd146, 8'd48, 1'b1, 1'b0};
2582: data_out = {8'd147, 8'd48, 1'b1, 1'b0};
2583: data_out = {8'd148, 8'd48, 1'b1, 1'b0};
2584: data_out = {8'd149, 8'd48, 1'b1, 1'b0};
2585: data_out = {8'd150, 8'd48, 1'b1, 1'b0};
2586: data_out = {8'd151, 8'd48, 1'b1, 1'b0};
2587: data_out = {8'd187, 8'd48, 1'b1, 1'b0};
2588: data_out = {8'd188, 8'd48, 1'b1, 1'b0};
2589: data_out = {8'd189, 8'd48, 1'b1, 1'b0};
2590: data_out = {8'd190, 8'd48, 1'b1, 1'b0};
2591: data_out = {8'd191, 8'd48, 1'b1, 1'b0};
2592: data_out = {8'd192, 8'd48, 1'b1, 1'b0};
2593: data_out = {8'd193, 8'd48, 1'b1, 1'b0};
2594: data_out = {8'd194, 8'd48, 1'b1, 1'b0};
2595: data_out = {8'd195, 8'd48, 1'b1, 1'b0};
2596: data_out = {8'd196, 8'd48, 1'b1, 1'b0};
2597: data_out = {8'd197, 8'd48, 1'b1, 1'b0};
2598: data_out = {8'd198, 8'd48, 1'b1, 1'b0};
2599: data_out = {8'd199, 8'd48, 1'b1, 1'b0};
2600: data_out = {8'd200, 8'd48, 1'b1, 1'b0};
2601: data_out = {8'd201, 8'd48, 1'b1, 1'b0};
2602: data_out = {8'd202, 8'd48, 1'b1, 1'b0};
2603: data_out = {8'd203, 8'd48, 1'b1, 1'b0};
2604: data_out = {8'd204, 8'd48, 1'b1, 1'b0};
2605: data_out = {8'd205, 8'd48, 1'b1, 1'b0};
2606: data_out = {8'd206, 8'd48, 1'b1, 1'b0};
2607: data_out = {8'd207, 8'd48, 1'b1, 1'b0};
2608: data_out = {8'd208, 8'd48, 1'b1, 1'b0};
2609: data_out = {8'd209, 8'd48, 1'b1, 1'b0};
2610: data_out = {8'd210, 8'd48, 1'b1, 1'b0};
2611: data_out = {8'd211, 8'd48, 1'b1, 1'b0};
2612: data_out = {8'd6, 8'd49, 1'b1, 1'b0};
2613: data_out = {8'd7, 8'd49, 1'b1, 1'b0};
2614: data_out = {8'd8, 8'd49, 1'b1, 1'b0};
2615: data_out = {8'd9, 8'd49, 1'b1, 1'b0};
2616: data_out = {8'd10, 8'd49, 1'b1, 1'b0};
2617: data_out = {8'd11, 8'd49, 1'b1, 1'b0};
2618: data_out = {8'd25, 8'd49, 1'b1, 1'b0};
2619: data_out = {8'd26, 8'd49, 1'b1, 1'b0};
2620: data_out = {8'd27, 8'd49, 1'b1, 1'b0};
2621: data_out = {8'd28, 8'd49, 1'b1, 1'b0};
2622: data_out = {8'd29, 8'd49, 1'b1, 1'b0};
2623: data_out = {8'd30, 8'd49, 1'b1, 1'b0};
2624: data_out = {8'd36, 8'd49, 1'b1, 1'b0};
2625: data_out = {8'd37, 8'd49, 1'b1, 1'b0};
2626: data_out = {8'd38, 8'd49, 1'b1, 1'b0};
2627: data_out = {8'd39, 8'd49, 1'b1, 1'b0};
2628: data_out = {8'd40, 8'd49, 1'b1, 1'b0};
2629: data_out = {8'd41, 8'd49, 1'b1, 1'b0};
2630: data_out = {8'd42, 8'd49, 1'b1, 1'b0};
2631: data_out = {8'd43, 8'd49, 1'b1, 1'b0};
2632: data_out = {8'd44, 8'd49, 1'b1, 1'b0};
2633: data_out = {8'd45, 8'd49, 1'b1, 1'b0};
2634: data_out = {8'd46, 8'd49, 1'b1, 1'b0};
2635: data_out = {8'd47, 8'd49, 1'b1, 1'b0};
2636: data_out = {8'd48, 8'd49, 1'b1, 1'b0};
2637: data_out = {8'd49, 8'd49, 1'b1, 1'b0};
2638: data_out = {8'd50, 8'd49, 1'b1, 1'b0};
2639: data_out = {8'd51, 8'd49, 1'b1, 1'b0};
2640: data_out = {8'd52, 8'd49, 1'b1, 1'b0};
2641: data_out = {8'd53, 8'd49, 1'b1, 1'b0};
2642: data_out = {8'd54, 8'd49, 1'b1, 1'b0};
2643: data_out = {8'd55, 8'd49, 1'b1, 1'b0};
2644: data_out = {8'd56, 8'd49, 1'b1, 1'b0};
2645: data_out = {8'd57, 8'd49, 1'b1, 1'b0};
2646: data_out = {8'd58, 8'd49, 1'b1, 1'b0};
2647: data_out = {8'd59, 8'd49, 1'b1, 1'b0};
2648: data_out = {8'd60, 8'd49, 1'b1, 1'b0};
2649: data_out = {8'd63, 8'd49, 1'b1, 1'b0};
2650: data_out = {8'd64, 8'd49, 1'b1, 1'b0};
2651: data_out = {8'd65, 8'd49, 1'b1, 1'b0};
2652: data_out = {8'd66, 8'd49, 1'b1, 1'b0};
2653: data_out = {8'd67, 8'd49, 1'b1, 1'b0};
2654: data_out = {8'd68, 8'd49, 1'b1, 1'b0};
2655: data_out = {8'd69, 8'd49, 1'b1, 1'b0};
2656: data_out = {8'd70, 8'd49, 1'b1, 1'b0};
2657: data_out = {8'd71, 8'd49, 1'b1, 1'b0};
2658: data_out = {8'd72, 8'd49, 1'b1, 1'b0};
2659: data_out = {8'd73, 8'd49, 1'b1, 1'b0};
2660: data_out = {8'd74, 8'd49, 1'b1, 1'b0};
2661: data_out = {8'd75, 8'd49, 1'b1, 1'b0};
2662: data_out = {8'd76, 8'd49, 1'b1, 1'b0};
2663: data_out = {8'd77, 8'd49, 1'b1, 1'b0};
2664: data_out = {8'd78, 8'd49, 1'b1, 1'b0};
2665: data_out = {8'd79, 8'd49, 1'b1, 1'b0};
2666: data_out = {8'd80, 8'd49, 1'b1, 1'b0};
2667: data_out = {8'd81, 8'd49, 1'b1, 1'b0};
2668: data_out = {8'd82, 8'd49, 1'b1, 1'b0};
2669: data_out = {8'd83, 8'd49, 1'b1, 1'b0};
2670: data_out = {8'd84, 8'd49, 1'b1, 1'b0};
2671: data_out = {8'd85, 8'd49, 1'b1, 1'b0};
2672: data_out = {8'd86, 8'd49, 1'b1, 1'b0};
2673: data_out = {8'd87, 8'd49, 1'b1, 1'b0};
2674: data_out = {8'd88, 8'd49, 1'b1, 1'b0};
2675: data_out = {8'd89, 8'd49, 1'b1, 1'b0};
2676: data_out = {8'd90, 8'd49, 1'b1, 1'b0};
2677: data_out = {8'd91, 8'd49, 1'b1, 1'b0};
2678: data_out = {8'd97, 8'd49, 1'b1, 1'b0};
2679: data_out = {8'd98, 8'd49, 1'b1, 1'b0};
2680: data_out = {8'd99, 8'd49, 1'b1, 1'b0};
2681: data_out = {8'd100, 8'd49, 1'b1, 1'b0};
2682: data_out = {8'd101, 8'd49, 1'b1, 1'b0};
2683: data_out = {8'd102, 8'd49, 1'b1, 1'b0};
2684: data_out = {8'd103, 8'd49, 1'b1, 1'b0};
2685: data_out = {8'd104, 8'd49, 1'b1, 1'b0};
2686: data_out = {8'd105, 8'd49, 1'b1, 1'b0};
2687: data_out = {8'd106, 8'd49, 1'b1, 1'b0};
2688: data_out = {8'd107, 8'd49, 1'b1, 1'b0};
2689: data_out = {8'd108, 8'd49, 1'b1, 1'b0};
2690: data_out = {8'd109, 8'd49, 1'b1, 1'b0};
2691: data_out = {8'd110, 8'd49, 1'b1, 1'b0};
2692: data_out = {8'd111, 8'd49, 1'b1, 1'b0};
2693: data_out = {8'd112, 8'd49, 1'b1, 1'b0};
2694: data_out = {8'd113, 8'd49, 1'b1, 1'b0};
2695: data_out = {8'd114, 8'd49, 1'b1, 1'b0};
2696: data_out = {8'd115, 8'd49, 1'b1, 1'b0};
2697: data_out = {8'd116, 8'd49, 1'b1, 1'b0};
2698: data_out = {8'd117, 8'd49, 1'b1, 1'b0};
2699: data_out = {8'd118, 8'd49, 1'b1, 1'b0};
2700: data_out = {8'd119, 8'd49, 1'b1, 1'b0};
2701: data_out = {8'd120, 8'd49, 1'b1, 1'b0};
2702: data_out = {8'd121, 8'd49, 1'b1, 1'b0};
2703: data_out = {8'd127, 8'd49, 1'b1, 1'b0};
2704: data_out = {8'd128, 8'd49, 1'b1, 1'b0};
2705: data_out = {8'd129, 8'd49, 1'b1, 1'b0};
2706: data_out = {8'd130, 8'd49, 1'b1, 1'b0};
2707: data_out = {8'd131, 8'd49, 1'b1, 1'b0};
2708: data_out = {8'd132, 8'd49, 1'b1, 1'b0};
2709: data_out = {8'd133, 8'd49, 1'b1, 1'b0};
2710: data_out = {8'd134, 8'd49, 1'b1, 1'b0};
2711: data_out = {8'd135, 8'd49, 1'b1, 1'b0};
2712: data_out = {8'd136, 8'd49, 1'b1, 1'b0};
2713: data_out = {8'd137, 8'd49, 1'b1, 1'b0};
2714: data_out = {8'd138, 8'd49, 1'b1, 1'b0};
2715: data_out = {8'd139, 8'd49, 1'b1, 1'b0};
2716: data_out = {8'd140, 8'd49, 1'b1, 1'b0};
2717: data_out = {8'd141, 8'd49, 1'b1, 1'b0};
2718: data_out = {8'd142, 8'd49, 1'b1, 1'b0};
2719: data_out = {8'd143, 8'd49, 1'b1, 1'b0};
2720: data_out = {8'd144, 8'd49, 1'b1, 1'b0};
2721: data_out = {8'd145, 8'd49, 1'b1, 1'b0};
2722: data_out = {8'd146, 8'd49, 1'b1, 1'b0};
2723: data_out = {8'd147, 8'd49, 1'b1, 1'b0};
2724: data_out = {8'd148, 8'd49, 1'b1, 1'b0};
2725: data_out = {8'd149, 8'd49, 1'b1, 1'b0};
2726: data_out = {8'd150, 8'd49, 1'b1, 1'b0};
2727: data_out = {8'd151, 8'd49, 1'b1, 1'b0};
2728: data_out = {8'd187, 8'd49, 1'b1, 1'b0};
2729: data_out = {8'd188, 8'd49, 1'b1, 1'b0};
2730: data_out = {8'd189, 8'd49, 1'b1, 1'b0};
2731: data_out = {8'd190, 8'd49, 1'b1, 1'b0};
2732: data_out = {8'd191, 8'd49, 1'b1, 1'b0};
2733: data_out = {8'd192, 8'd49, 1'b1, 1'b0};
2734: data_out = {8'd193, 8'd49, 1'b1, 1'b0};
2735: data_out = {8'd194, 8'd49, 1'b1, 1'b0};
2736: data_out = {8'd195, 8'd49, 1'b1, 1'b0};
2737: data_out = {8'd196, 8'd49, 1'b1, 1'b0};
2738: data_out = {8'd197, 8'd49, 1'b1, 1'b0};
2739: data_out = {8'd198, 8'd49, 1'b1, 1'b0};
2740: data_out = {8'd199, 8'd49, 1'b1, 1'b0};
2741: data_out = {8'd200, 8'd49, 1'b1, 1'b0};
2742: data_out = {8'd201, 8'd49, 1'b1, 1'b0};
2743: data_out = {8'd202, 8'd49, 1'b1, 1'b0};
2744: data_out = {8'd203, 8'd49, 1'b1, 1'b0};
2745: data_out = {8'd204, 8'd49, 1'b1, 1'b0};
2746: data_out = {8'd205, 8'd49, 1'b1, 1'b0};
2747: data_out = {8'd206, 8'd49, 1'b1, 1'b0};
2748: data_out = {8'd207, 8'd49, 1'b1, 1'b0};
2749: data_out = {8'd208, 8'd49, 1'b1, 1'b0};
2750: data_out = {8'd209, 8'd49, 1'b1, 1'b0};
2751: data_out = {8'd210, 8'd49, 1'b1, 1'b0};
2752: data_out = {8'd211, 8'd49, 1'b1, 1'b0};
2753: data_out = {8'd6, 8'd50, 1'b1, 1'b0};
2754: data_out = {8'd7, 8'd50, 1'b1, 1'b0};
2755: data_out = {8'd8, 8'd50, 1'b1, 1'b0};
2756: data_out = {8'd9, 8'd50, 1'b1, 1'b0};
2757: data_out = {8'd10, 8'd50, 1'b1, 1'b0};
2758: data_out = {8'd11, 8'd50, 1'b1, 1'b0};
2759: data_out = {8'd25, 8'd50, 1'b1, 1'b0};
2760: data_out = {8'd26, 8'd50, 1'b1, 1'b0};
2761: data_out = {8'd27, 8'd50, 1'b1, 1'b0};
2762: data_out = {8'd28, 8'd50, 1'b1, 1'b0};
2763: data_out = {8'd29, 8'd50, 1'b1, 1'b0};
2764: data_out = {8'd30, 8'd50, 1'b1, 1'b0};
2765: data_out = {8'd36, 8'd50, 1'b1, 1'b0};
2766: data_out = {8'd37, 8'd50, 1'b1, 1'b0};
2767: data_out = {8'd38, 8'd50, 1'b1, 1'b0};
2768: data_out = {8'd39, 8'd50, 1'b1, 1'b0};
2769: data_out = {8'd40, 8'd50, 1'b1, 1'b0};
2770: data_out = {8'd41, 8'd50, 1'b1, 1'b0};
2771: data_out = {8'd42, 8'd50, 1'b1, 1'b0};
2772: data_out = {8'd43, 8'd50, 1'b1, 1'b0};
2773: data_out = {8'd44, 8'd50, 1'b1, 1'b0};
2774: data_out = {8'd45, 8'd50, 1'b1, 1'b0};
2775: data_out = {8'd46, 8'd50, 1'b1, 1'b0};
2776: data_out = {8'd47, 8'd50, 1'b1, 1'b0};
2777: data_out = {8'd48, 8'd50, 1'b1, 1'b0};
2778: data_out = {8'd49, 8'd50, 1'b1, 1'b0};
2779: data_out = {8'd50, 8'd50, 1'b1, 1'b0};
2780: data_out = {8'd51, 8'd50, 1'b1, 1'b0};
2781: data_out = {8'd52, 8'd50, 1'b1, 1'b0};
2782: data_out = {8'd53, 8'd50, 1'b1, 1'b0};
2783: data_out = {8'd54, 8'd50, 1'b1, 1'b0};
2784: data_out = {8'd55, 8'd50, 1'b1, 1'b0};
2785: data_out = {8'd56, 8'd50, 1'b1, 1'b0};
2786: data_out = {8'd57, 8'd50, 1'b1, 1'b0};
2787: data_out = {8'd58, 8'd50, 1'b1, 1'b0};
2788: data_out = {8'd59, 8'd50, 1'b1, 1'b0};
2789: data_out = {8'd60, 8'd50, 1'b1, 1'b0};
2790: data_out = {8'd63, 8'd50, 1'b1, 1'b0};
2791: data_out = {8'd64, 8'd50, 1'b1, 1'b0};
2792: data_out = {8'd65, 8'd50, 1'b1, 1'b0};
2793: data_out = {8'd66, 8'd50, 1'b1, 1'b0};
2794: data_out = {8'd67, 8'd50, 1'b1, 1'b0};
2795: data_out = {8'd68, 8'd50, 1'b1, 1'b0};
2796: data_out = {8'd69, 8'd50, 1'b1, 1'b0};
2797: data_out = {8'd70, 8'd50, 1'b1, 1'b0};
2798: data_out = {8'd71, 8'd50, 1'b1, 1'b0};
2799: data_out = {8'd72, 8'd50, 1'b1, 1'b0};
2800: data_out = {8'd73, 8'd50, 1'b1, 1'b0};
2801: data_out = {8'd74, 8'd50, 1'b1, 1'b0};
2802: data_out = {8'd75, 8'd50, 1'b1, 1'b0};
2803: data_out = {8'd76, 8'd50, 1'b1, 1'b0};
2804: data_out = {8'd77, 8'd50, 1'b1, 1'b0};
2805: data_out = {8'd78, 8'd50, 1'b1, 1'b0};
2806: data_out = {8'd79, 8'd50, 1'b1, 1'b0};
2807: data_out = {8'd80, 8'd50, 1'b1, 1'b0};
2808: data_out = {8'd81, 8'd50, 1'b1, 1'b0};
2809: data_out = {8'd82, 8'd50, 1'b1, 1'b0};
2810: data_out = {8'd83, 8'd50, 1'b1, 1'b0};
2811: data_out = {8'd84, 8'd50, 1'b1, 1'b0};
2812: data_out = {8'd85, 8'd50, 1'b1, 1'b0};
2813: data_out = {8'd86, 8'd50, 1'b1, 1'b0};
2814: data_out = {8'd87, 8'd50, 1'b1, 1'b0};
2815: data_out = {8'd88, 8'd50, 1'b1, 1'b0};
2816: data_out = {8'd89, 8'd50, 1'b1, 1'b0};
2817: data_out = {8'd90, 8'd50, 1'b1, 1'b0};
2818: data_out = {8'd91, 8'd50, 1'b1, 1'b0};
2819: data_out = {8'd97, 8'd50, 1'b1, 1'b0};
2820: data_out = {8'd98, 8'd50, 1'b1, 1'b0};
2821: data_out = {8'd99, 8'd50, 1'b1, 1'b0};
2822: data_out = {8'd100, 8'd50, 1'b1, 1'b0};
2823: data_out = {8'd101, 8'd50, 1'b1, 1'b0};
2824: data_out = {8'd102, 8'd50, 1'b1, 1'b0};
2825: data_out = {8'd103, 8'd50, 1'b1, 1'b0};
2826: data_out = {8'd104, 8'd50, 1'b1, 1'b0};
2827: data_out = {8'd105, 8'd50, 1'b1, 1'b0};
2828: data_out = {8'd106, 8'd50, 1'b1, 1'b0};
2829: data_out = {8'd107, 8'd50, 1'b1, 1'b0};
2830: data_out = {8'd108, 8'd50, 1'b1, 1'b0};
2831: data_out = {8'd109, 8'd50, 1'b1, 1'b0};
2832: data_out = {8'd110, 8'd50, 1'b1, 1'b0};
2833: data_out = {8'd111, 8'd50, 1'b1, 1'b0};
2834: data_out = {8'd112, 8'd50, 1'b1, 1'b0};
2835: data_out = {8'd113, 8'd50, 1'b1, 1'b0};
2836: data_out = {8'd114, 8'd50, 1'b1, 1'b0};
2837: data_out = {8'd115, 8'd50, 1'b1, 1'b0};
2838: data_out = {8'd116, 8'd50, 1'b1, 1'b0};
2839: data_out = {8'd117, 8'd50, 1'b1, 1'b0};
2840: data_out = {8'd118, 8'd50, 1'b1, 1'b0};
2841: data_out = {8'd119, 8'd50, 1'b1, 1'b0};
2842: data_out = {8'd120, 8'd50, 1'b1, 1'b0};
2843: data_out = {8'd121, 8'd50, 1'b1, 1'b0};
2844: data_out = {8'd127, 8'd50, 1'b1, 1'b0};
2845: data_out = {8'd128, 8'd50, 1'b1, 1'b0};
2846: data_out = {8'd129, 8'd50, 1'b1, 1'b0};
2847: data_out = {8'd130, 8'd50, 1'b1, 1'b0};
2848: data_out = {8'd131, 8'd50, 1'b1, 1'b0};
2849: data_out = {8'd132, 8'd50, 1'b1, 1'b0};
2850: data_out = {8'd133, 8'd50, 1'b1, 1'b0};
2851: data_out = {8'd134, 8'd50, 1'b1, 1'b0};
2852: data_out = {8'd135, 8'd50, 1'b1, 1'b0};
2853: data_out = {8'd136, 8'd50, 1'b1, 1'b0};
2854: data_out = {8'd137, 8'd50, 1'b1, 1'b0};
2855: data_out = {8'd138, 8'd50, 1'b1, 1'b0};
2856: data_out = {8'd139, 8'd50, 1'b1, 1'b0};
2857: data_out = {8'd140, 8'd50, 1'b1, 1'b0};
2858: data_out = {8'd141, 8'd50, 1'b1, 1'b0};
2859: data_out = {8'd142, 8'd50, 1'b1, 1'b0};
2860: data_out = {8'd143, 8'd50, 1'b1, 1'b0};
2861: data_out = {8'd144, 8'd50, 1'b1, 1'b0};
2862: data_out = {8'd145, 8'd50, 1'b1, 1'b0};
2863: data_out = {8'd146, 8'd50, 1'b1, 1'b0};
2864: data_out = {8'd147, 8'd50, 1'b1, 1'b0};
2865: data_out = {8'd148, 8'd50, 1'b1, 1'b0};
2866: data_out = {8'd149, 8'd50, 1'b1, 1'b0};
2867: data_out = {8'd150, 8'd50, 1'b1, 1'b0};
2868: data_out = {8'd151, 8'd50, 1'b1, 1'b0};
2869: data_out = {8'd187, 8'd50, 1'b1, 1'b0};
2870: data_out = {8'd188, 8'd50, 1'b1, 1'b0};
2871: data_out = {8'd189, 8'd50, 1'b1, 1'b0};
2872: data_out = {8'd190, 8'd50, 1'b1, 1'b0};
2873: data_out = {8'd191, 8'd50, 1'b1, 1'b0};
2874: data_out = {8'd192, 8'd50, 1'b1, 1'b0};
2875: data_out = {8'd193, 8'd50, 1'b1, 1'b0};
2876: data_out = {8'd194, 8'd50, 1'b1, 1'b0};
2877: data_out = {8'd195, 8'd50, 1'b1, 1'b0};
2878: data_out = {8'd196, 8'd50, 1'b1, 1'b0};
2879: data_out = {8'd197, 8'd50, 1'b1, 1'b0};
2880: data_out = {8'd198, 8'd50, 1'b1, 1'b0};
2881: data_out = {8'd199, 8'd50, 1'b1, 1'b0};
2882: data_out = {8'd200, 8'd50, 1'b1, 1'b0};
2883: data_out = {8'd201, 8'd50, 1'b1, 1'b0};
2884: data_out = {8'd202, 8'd50, 1'b1, 1'b0};
2885: data_out = {8'd203, 8'd50, 1'b1, 1'b0};
2886: data_out = {8'd204, 8'd50, 1'b1, 1'b0};
2887: data_out = {8'd205, 8'd50, 1'b1, 1'b0};
2888: data_out = {8'd206, 8'd50, 1'b1, 1'b0};
2889: data_out = {8'd207, 8'd50, 1'b1, 1'b0};
2890: data_out = {8'd208, 8'd50, 1'b1, 1'b0};
2891: data_out = {8'd209, 8'd50, 1'b1, 1'b0};
2892: data_out = {8'd210, 8'd50, 1'b1, 1'b0};
2893: data_out = {8'd211, 8'd50, 1'b1, 1'b0};
2894: data_out = {8'd6, 8'd51, 1'b1, 1'b0};
2895: data_out = {8'd7, 8'd51, 1'b1, 1'b0};
2896: data_out = {8'd8, 8'd51, 1'b1, 1'b0};
2897: data_out = {8'd9, 8'd51, 1'b1, 1'b0};
2898: data_out = {8'd10, 8'd51, 1'b1, 1'b0};
2899: data_out = {8'd11, 8'd51, 1'b1, 1'b0};
2900: data_out = {8'd25, 8'd51, 1'b1, 1'b0};
2901: data_out = {8'd26, 8'd51, 1'b1, 1'b0};
2902: data_out = {8'd27, 8'd51, 1'b1, 1'b0};
2903: data_out = {8'd28, 8'd51, 1'b1, 1'b0};
2904: data_out = {8'd29, 8'd51, 1'b1, 1'b0};
2905: data_out = {8'd30, 8'd51, 1'b1, 1'b0};
2906: data_out = {8'd37, 8'd51, 1'b1, 1'b0};
2907: data_out = {8'd38, 8'd51, 1'b1, 1'b0};
2908: data_out = {8'd39, 8'd51, 1'b1, 1'b0};
2909: data_out = {8'd40, 8'd51, 1'b1, 1'b0};
2910: data_out = {8'd41, 8'd51, 1'b1, 1'b0};
2911: data_out = {8'd42, 8'd51, 1'b1, 1'b0};
2912: data_out = {8'd43, 8'd51, 1'b1, 1'b0};
2913: data_out = {8'd44, 8'd51, 1'b1, 1'b0};
2914: data_out = {8'd45, 8'd51, 1'b1, 1'b0};
2915: data_out = {8'd46, 8'd51, 1'b1, 1'b0};
2916: data_out = {8'd47, 8'd51, 1'b1, 1'b0};
2917: data_out = {8'd48, 8'd51, 1'b1, 1'b0};
2918: data_out = {8'd49, 8'd51, 1'b1, 1'b0};
2919: data_out = {8'd50, 8'd51, 1'b1, 1'b0};
2920: data_out = {8'd51, 8'd51, 1'b1, 1'b0};
2921: data_out = {8'd52, 8'd51, 1'b1, 1'b0};
2922: data_out = {8'd53, 8'd51, 1'b1, 1'b0};
2923: data_out = {8'd54, 8'd51, 1'b1, 1'b0};
2924: data_out = {8'd55, 8'd51, 1'b1, 1'b0};
2925: data_out = {8'd56, 8'd51, 1'b1, 1'b0};
2926: data_out = {8'd57, 8'd51, 1'b1, 1'b0};
2927: data_out = {8'd58, 8'd51, 1'b1, 1'b0};
2928: data_out = {8'd59, 8'd51, 1'b1, 1'b0};
2929: data_out = {8'd63, 8'd51, 1'b1, 1'b0};
2930: data_out = {8'd64, 8'd51, 1'b1, 1'b0};
2931: data_out = {8'd65, 8'd51, 1'b1, 1'b0};
2932: data_out = {8'd66, 8'd51, 1'b1, 1'b0};
2933: data_out = {8'd67, 8'd51, 1'b1, 1'b0};
2934: data_out = {8'd68, 8'd51, 1'b1, 1'b0};
2935: data_out = {8'd69, 8'd51, 1'b1, 1'b0};
2936: data_out = {8'd70, 8'd51, 1'b1, 1'b0};
2937: data_out = {8'd71, 8'd51, 1'b1, 1'b0};
2938: data_out = {8'd72, 8'd51, 1'b1, 1'b0};
2939: data_out = {8'd73, 8'd51, 1'b1, 1'b0};
2940: data_out = {8'd74, 8'd51, 1'b1, 1'b0};
2941: data_out = {8'd75, 8'd51, 1'b1, 1'b0};
2942: data_out = {8'd76, 8'd51, 1'b1, 1'b0};
2943: data_out = {8'd77, 8'd51, 1'b1, 1'b0};
2944: data_out = {8'd78, 8'd51, 1'b1, 1'b0};
2945: data_out = {8'd79, 8'd51, 1'b1, 1'b0};
2946: data_out = {8'd80, 8'd51, 1'b1, 1'b0};
2947: data_out = {8'd81, 8'd51, 1'b1, 1'b0};
2948: data_out = {8'd82, 8'd51, 1'b1, 1'b0};
2949: data_out = {8'd83, 8'd51, 1'b1, 1'b0};
2950: data_out = {8'd84, 8'd51, 1'b1, 1'b0};
2951: data_out = {8'd85, 8'd51, 1'b1, 1'b0};
2952: data_out = {8'd86, 8'd51, 1'b1, 1'b0};
2953: data_out = {8'd87, 8'd51, 1'b1, 1'b0};
2954: data_out = {8'd88, 8'd51, 1'b1, 1'b0};
2955: data_out = {8'd89, 8'd51, 1'b1, 1'b0};
2956: data_out = {8'd90, 8'd51, 1'b1, 1'b0};
2957: data_out = {8'd91, 8'd51, 1'b1, 1'b0};
2958: data_out = {8'd98, 8'd51, 1'b1, 1'b0};
2959: data_out = {8'd99, 8'd51, 1'b1, 1'b0};
2960: data_out = {8'd100, 8'd51, 1'b1, 1'b0};
2961: data_out = {8'd101, 8'd51, 1'b1, 1'b0};
2962: data_out = {8'd102, 8'd51, 1'b1, 1'b0};
2963: data_out = {8'd103, 8'd51, 1'b1, 1'b0};
2964: data_out = {8'd104, 8'd51, 1'b1, 1'b0};
2965: data_out = {8'd105, 8'd51, 1'b1, 1'b0};
2966: data_out = {8'd106, 8'd51, 1'b1, 1'b0};
2967: data_out = {8'd107, 8'd51, 1'b1, 1'b0};
2968: data_out = {8'd108, 8'd51, 1'b1, 1'b0};
2969: data_out = {8'd109, 8'd51, 1'b1, 1'b0};
2970: data_out = {8'd110, 8'd51, 1'b1, 1'b0};
2971: data_out = {8'd111, 8'd51, 1'b1, 1'b0};
2972: data_out = {8'd112, 8'd51, 1'b1, 1'b0};
2973: data_out = {8'd113, 8'd51, 1'b1, 1'b0};
2974: data_out = {8'd114, 8'd51, 1'b1, 1'b0};
2975: data_out = {8'd115, 8'd51, 1'b1, 1'b0};
2976: data_out = {8'd116, 8'd51, 1'b1, 1'b0};
2977: data_out = {8'd117, 8'd51, 1'b1, 1'b0};
2978: data_out = {8'd118, 8'd51, 1'b1, 1'b0};
2979: data_out = {8'd119, 8'd51, 1'b1, 1'b0};
2980: data_out = {8'd120, 8'd51, 1'b1, 1'b0};
2981: data_out = {8'd128, 8'd51, 1'b1, 1'b0};
2982: data_out = {8'd129, 8'd51, 1'b1, 1'b0};
2983: data_out = {8'd130, 8'd51, 1'b1, 1'b0};
2984: data_out = {8'd131, 8'd51, 1'b1, 1'b0};
2985: data_out = {8'd132, 8'd51, 1'b1, 1'b0};
2986: data_out = {8'd133, 8'd51, 1'b1, 1'b0};
2987: data_out = {8'd134, 8'd51, 1'b1, 1'b0};
2988: data_out = {8'd135, 8'd51, 1'b1, 1'b0};
2989: data_out = {8'd136, 8'd51, 1'b1, 1'b0};
2990: data_out = {8'd137, 8'd51, 1'b1, 1'b0};
2991: data_out = {8'd138, 8'd51, 1'b1, 1'b0};
2992: data_out = {8'd139, 8'd51, 1'b1, 1'b0};
2993: data_out = {8'd140, 8'd51, 1'b1, 1'b0};
2994: data_out = {8'd141, 8'd51, 1'b1, 1'b0};
2995: data_out = {8'd142, 8'd51, 1'b1, 1'b0};
2996: data_out = {8'd143, 8'd51, 1'b1, 1'b0};
2997: data_out = {8'd144, 8'd51, 1'b1, 1'b0};
2998: data_out = {8'd145, 8'd51, 1'b1, 1'b0};
2999: data_out = {8'd146, 8'd51, 1'b1, 1'b0};
3000: data_out = {8'd147, 8'd51, 1'b1, 1'b0};
3001: data_out = {8'd148, 8'd51, 1'b1, 1'b0};
3002: data_out = {8'd149, 8'd51, 1'b1, 1'b0};
3003: data_out = {8'd150, 8'd51, 1'b1, 1'b0};
3004: data_out = {8'd188, 8'd51, 1'b1, 1'b0};
3005: data_out = {8'd189, 8'd51, 1'b1, 1'b0};
3006: data_out = {8'd190, 8'd51, 1'b1, 1'b0};
3007: data_out = {8'd191, 8'd51, 1'b1, 1'b0};
3008: data_out = {8'd192, 8'd51, 1'b1, 1'b0};
3009: data_out = {8'd193, 8'd51, 1'b1, 1'b0};
3010: data_out = {8'd194, 8'd51, 1'b1, 1'b0};
3011: data_out = {8'd195, 8'd51, 1'b1, 1'b0};
3012: data_out = {8'd196, 8'd51, 1'b1, 1'b0};
3013: data_out = {8'd197, 8'd51, 1'b1, 1'b0};
3014: data_out = {8'd198, 8'd51, 1'b1, 1'b0};
3015: data_out = {8'd199, 8'd51, 1'b1, 1'b0};
3016: data_out = {8'd200, 8'd51, 1'b1, 1'b0};
3017: data_out = {8'd201, 8'd51, 1'b1, 1'b0};
3018: data_out = {8'd202, 8'd51, 1'b1, 1'b0};
3019: data_out = {8'd203, 8'd51, 1'b1, 1'b0};
3020: data_out = {8'd204, 8'd51, 1'b1, 1'b0};
3021: data_out = {8'd205, 8'd51, 1'b1, 1'b0};
3022: data_out = {8'd206, 8'd51, 1'b1, 1'b0};
3023: data_out = {8'd207, 8'd51, 1'b1, 1'b0};
3024: data_out = {8'd208, 8'd51, 1'b1, 1'b0};
3025: data_out = {8'd209, 8'd51, 1'b1, 1'b0};
3026: data_out = {8'd210, 8'd51, 1'b1, 1'b0};
3027: data_out = {8'd6, 8'd52, 1'b1, 1'b0};
3028: data_out = {8'd7, 8'd52, 1'b1, 1'b0};
3029: data_out = {8'd8, 8'd52, 1'b1, 1'b0};
3030: data_out = {8'd9, 8'd52, 1'b1, 1'b0};
3031: data_out = {8'd10, 8'd52, 1'b1, 1'b0};
3032: data_out = {8'd11, 8'd52, 1'b1, 1'b0};
3033: data_out = {8'd25, 8'd52, 1'b1, 1'b0};
3034: data_out = {8'd26, 8'd52, 1'b1, 1'b0};
3035: data_out = {8'd27, 8'd52, 1'b1, 1'b0};
3036: data_out = {8'd28, 8'd52, 1'b1, 1'b0};
3037: data_out = {8'd29, 8'd52, 1'b1, 1'b0};
3038: data_out = {8'd30, 8'd52, 1'b1, 1'b0};
3039: data_out = {8'd38, 8'd52, 1'b1, 1'b0};
3040: data_out = {8'd39, 8'd52, 1'b1, 1'b0};
3041: data_out = {8'd40, 8'd52, 1'b1, 1'b0};
3042: data_out = {8'd41, 8'd52, 1'b1, 1'b0};
3043: data_out = {8'd42, 8'd52, 1'b1, 1'b0};
3044: data_out = {8'd43, 8'd52, 1'b1, 1'b0};
3045: data_out = {8'd44, 8'd52, 1'b1, 1'b0};
3046: data_out = {8'd45, 8'd52, 1'b1, 1'b0};
3047: data_out = {8'd46, 8'd52, 1'b1, 1'b0};
3048: data_out = {8'd47, 8'd52, 1'b1, 1'b0};
3049: data_out = {8'd48, 8'd52, 1'b1, 1'b0};
3050: data_out = {8'd49, 8'd52, 1'b1, 1'b0};
3051: data_out = {8'd50, 8'd52, 1'b1, 1'b0};
3052: data_out = {8'd51, 8'd52, 1'b1, 1'b0};
3053: data_out = {8'd52, 8'd52, 1'b1, 1'b0};
3054: data_out = {8'd53, 8'd52, 1'b1, 1'b0};
3055: data_out = {8'd54, 8'd52, 1'b1, 1'b0};
3056: data_out = {8'd55, 8'd52, 1'b1, 1'b0};
3057: data_out = {8'd56, 8'd52, 1'b1, 1'b0};
3058: data_out = {8'd57, 8'd52, 1'b1, 1'b0};
3059: data_out = {8'd58, 8'd52, 1'b1, 1'b0};
3060: data_out = {8'd63, 8'd52, 1'b1, 1'b0};
3061: data_out = {8'd64, 8'd52, 1'b1, 1'b0};
3062: data_out = {8'd65, 8'd52, 1'b1, 1'b0};
3063: data_out = {8'd66, 8'd52, 1'b1, 1'b0};
3064: data_out = {8'd67, 8'd52, 1'b1, 1'b0};
3065: data_out = {8'd68, 8'd52, 1'b1, 1'b0};
3066: data_out = {8'd69, 8'd52, 1'b1, 1'b0};
3067: data_out = {8'd70, 8'd52, 1'b1, 1'b0};
3068: data_out = {8'd71, 8'd52, 1'b1, 1'b0};
3069: data_out = {8'd72, 8'd52, 1'b1, 1'b0};
3070: data_out = {8'd73, 8'd52, 1'b1, 1'b0};
3071: data_out = {8'd74, 8'd52, 1'b1, 1'b0};
3072: data_out = {8'd75, 8'd52, 1'b1, 1'b0};
3073: data_out = {8'd76, 8'd52, 1'b1, 1'b0};
3074: data_out = {8'd77, 8'd52, 1'b1, 1'b0};
3075: data_out = {8'd78, 8'd52, 1'b1, 1'b0};
3076: data_out = {8'd79, 8'd52, 1'b1, 1'b0};
3077: data_out = {8'd80, 8'd52, 1'b1, 1'b0};
3078: data_out = {8'd81, 8'd52, 1'b1, 1'b0};
3079: data_out = {8'd82, 8'd52, 1'b1, 1'b0};
3080: data_out = {8'd83, 8'd52, 1'b1, 1'b0};
3081: data_out = {8'd84, 8'd52, 1'b1, 1'b0};
3082: data_out = {8'd85, 8'd52, 1'b1, 1'b0};
3083: data_out = {8'd86, 8'd52, 1'b1, 1'b0};
3084: data_out = {8'd87, 8'd52, 1'b1, 1'b0};
3085: data_out = {8'd88, 8'd52, 1'b1, 1'b0};
3086: data_out = {8'd89, 8'd52, 1'b1, 1'b0};
3087: data_out = {8'd90, 8'd52, 1'b1, 1'b0};
3088: data_out = {8'd91, 8'd52, 1'b1, 1'b0};
3089: data_out = {8'd99, 8'd52, 1'b1, 1'b0};
3090: data_out = {8'd100, 8'd52, 1'b1, 1'b0};
3091: data_out = {8'd101, 8'd52, 1'b1, 1'b0};
3092: data_out = {8'd102, 8'd52, 1'b1, 1'b0};
3093: data_out = {8'd103, 8'd52, 1'b1, 1'b0};
3094: data_out = {8'd104, 8'd52, 1'b1, 1'b0};
3095: data_out = {8'd105, 8'd52, 1'b1, 1'b0};
3096: data_out = {8'd106, 8'd52, 1'b1, 1'b0};
3097: data_out = {8'd107, 8'd52, 1'b1, 1'b0};
3098: data_out = {8'd108, 8'd52, 1'b1, 1'b0};
3099: data_out = {8'd109, 8'd52, 1'b1, 1'b0};
3100: data_out = {8'd110, 8'd52, 1'b1, 1'b0};
3101: data_out = {8'd111, 8'd52, 1'b1, 1'b0};
3102: data_out = {8'd112, 8'd52, 1'b1, 1'b0};
3103: data_out = {8'd113, 8'd52, 1'b1, 1'b0};
3104: data_out = {8'd114, 8'd52, 1'b1, 1'b0};
3105: data_out = {8'd115, 8'd52, 1'b1, 1'b0};
3106: data_out = {8'd116, 8'd52, 1'b1, 1'b0};
3107: data_out = {8'd117, 8'd52, 1'b1, 1'b0};
3108: data_out = {8'd118, 8'd52, 1'b1, 1'b0};
3109: data_out = {8'd119, 8'd52, 1'b1, 1'b0};
3110: data_out = {8'd129, 8'd52, 1'b1, 1'b0};
3111: data_out = {8'd130, 8'd52, 1'b1, 1'b0};
3112: data_out = {8'd131, 8'd52, 1'b1, 1'b0};
3113: data_out = {8'd132, 8'd52, 1'b1, 1'b0};
3114: data_out = {8'd133, 8'd52, 1'b1, 1'b0};
3115: data_out = {8'd134, 8'd52, 1'b1, 1'b0};
3116: data_out = {8'd135, 8'd52, 1'b1, 1'b0};
3117: data_out = {8'd136, 8'd52, 1'b1, 1'b0};
3118: data_out = {8'd137, 8'd52, 1'b1, 1'b0};
3119: data_out = {8'd138, 8'd52, 1'b1, 1'b0};
3120: data_out = {8'd139, 8'd52, 1'b1, 1'b0};
3121: data_out = {8'd140, 8'd52, 1'b1, 1'b0};
3122: data_out = {8'd141, 8'd52, 1'b1, 1'b0};
3123: data_out = {8'd142, 8'd52, 1'b1, 1'b0};
3124: data_out = {8'd143, 8'd52, 1'b1, 1'b0};
3125: data_out = {8'd144, 8'd52, 1'b1, 1'b0};
3126: data_out = {8'd145, 8'd52, 1'b1, 1'b0};
3127: data_out = {8'd146, 8'd52, 1'b1, 1'b0};
3128: data_out = {8'd147, 8'd52, 1'b1, 1'b0};
3129: data_out = {8'd148, 8'd52, 1'b1, 1'b0};
3130: data_out = {8'd149, 8'd52, 1'b1, 1'b0};
3131: data_out = {8'd189, 8'd52, 1'b1, 1'b0};
3132: data_out = {8'd190, 8'd52, 1'b1, 1'b0};
3133: data_out = {8'd191, 8'd52, 1'b1, 1'b0};
3134: data_out = {8'd192, 8'd52, 1'b1, 1'b0};
3135: data_out = {8'd193, 8'd52, 1'b1, 1'b0};
3136: data_out = {8'd194, 8'd52, 1'b1, 1'b0};
3137: data_out = {8'd195, 8'd52, 1'b1, 1'b0};
3138: data_out = {8'd196, 8'd52, 1'b1, 1'b0};
3139: data_out = {8'd197, 8'd52, 1'b1, 1'b0};
3140: data_out = {8'd198, 8'd52, 1'b1, 1'b0};
3141: data_out = {8'd199, 8'd52, 1'b1, 1'b0};
3142: data_out = {8'd200, 8'd52, 1'b1, 1'b0};
3143: data_out = {8'd201, 8'd52, 1'b1, 1'b0};
3144: data_out = {8'd202, 8'd52, 1'b1, 1'b0};
3145: data_out = {8'd203, 8'd52, 1'b1, 1'b0};
3146: data_out = {8'd204, 8'd52, 1'b1, 1'b0};
3147: data_out = {8'd205, 8'd52, 1'b1, 1'b0};
3148: data_out = {8'd206, 8'd52, 1'b1, 1'b0};
3149: data_out = {8'd207, 8'd52, 1'b1, 1'b0};
3150: data_out = {8'd208, 8'd52, 1'b1, 1'b0};
3151: data_out = {8'd209, 8'd52, 1'b1, 1'b0};
3152: data_out = {8'd70, 8'd74, 1'b1, 1'b0};
3153: data_out = {8'd157, 8'd74, 1'b1, 1'b0};
3154: data_out = {8'd70, 8'd75, 1'b1, 1'b0};
3155: data_out = {8'd100, 8'd75, 1'b1, 1'b0};
3156: data_out = {8'd6, 8'd76, 1'b1, 1'b0};
3157: data_out = {8'd7, 8'd76, 1'b1, 1'b0};
3158: data_out = {8'd8, 8'd76, 1'b1, 1'b0};
3159: data_out = {8'd9, 8'd76, 1'b1, 1'b0};
3160: data_out = {8'd10, 8'd76, 1'b1, 1'b0};
3161: data_out = {8'd13, 8'd76, 1'b1, 1'b0};
3162: data_out = {8'd14, 8'd76, 1'b1, 1'b0};
3163: data_out = {8'd15, 8'd76, 1'b1, 1'b0};
3164: data_out = {8'd16, 8'd76, 1'b1, 1'b0};
3165: data_out = {8'd17, 8'd76, 1'b1, 1'b0};
3166: data_out = {8'd26, 8'd76, 1'b1, 1'b0};
3167: data_out = {8'd27, 8'd76, 1'b1, 1'b0};
3168: data_out = {8'd28, 8'd76, 1'b1, 1'b0};
3169: data_out = {8'd29, 8'd76, 1'b1, 1'b0};
3170: data_out = {8'd30, 8'd76, 1'b1, 1'b0};
3171: data_out = {8'd39, 8'd76, 1'b1, 1'b0};
3172: data_out = {8'd40, 8'd76, 1'b1, 1'b0};
3173: data_out = {8'd41, 8'd76, 1'b1, 1'b0};
3174: data_out = {8'd42, 8'd76, 1'b1, 1'b0};
3175: data_out = {8'd43, 8'd76, 1'b1, 1'b0};
3176: data_out = {8'd46, 8'd76, 1'b1, 1'b0};
3177: data_out = {8'd47, 8'd76, 1'b1, 1'b0};
3178: data_out = {8'd48, 8'd76, 1'b1, 1'b0};
3179: data_out = {8'd49, 8'd76, 1'b1, 1'b0};
3180: data_out = {8'd50, 8'd76, 1'b1, 1'b0};
3181: data_out = {8'd54, 8'd76, 1'b1, 1'b0};
3182: data_out = {8'd55, 8'd76, 1'b1, 1'b0};
3183: data_out = {8'd56, 8'd76, 1'b1, 1'b0};
3184: data_out = {8'd59, 8'd76, 1'b1, 1'b0};
3185: data_out = {8'd60, 8'd76, 1'b1, 1'b0};
3186: data_out = {8'd61, 8'd76, 1'b1, 1'b0};
3187: data_out = {8'd62, 8'd76, 1'b1, 1'b0};
3188: data_out = {8'd63, 8'd76, 1'b1, 1'b0};
3189: data_out = {8'd66, 8'd76, 1'b1, 1'b0};
3190: data_out = {8'd67, 8'd76, 1'b1, 1'b0};
3191: data_out = {8'd68, 8'd76, 1'b1, 1'b0};
3192: data_out = {8'd69, 8'd76, 1'b1, 1'b0};
3193: data_out = {8'd70, 8'd76, 1'b1, 1'b0};
3194: data_out = {8'd79, 8'd76, 1'b1, 1'b0};
3195: data_out = {8'd80, 8'd76, 1'b1, 1'b0};
3196: data_out = {8'd81, 8'd76, 1'b1, 1'b0};
3197: data_out = {8'd82, 8'd76, 1'b1, 1'b0};
3198: data_out = {8'd83, 8'd76, 1'b1, 1'b0};
3199: data_out = {8'd86, 8'd76, 1'b1, 1'b0};
3200: data_out = {8'd90, 8'd76, 1'b1, 1'b0};
3201: data_out = {8'd93, 8'd76, 1'b1, 1'b0};
3202: data_out = {8'd94, 8'd76, 1'b1, 1'b0};
3203: data_out = {8'd95, 8'd76, 1'b1, 1'b0};
3204: data_out = {8'd96, 8'd76, 1'b1, 1'b0};
3205: data_out = {8'd97, 8'd76, 1'b1, 1'b0};
3206: data_out = {8'd99, 8'd76, 1'b1, 1'b0};
3207: data_out = {8'd100, 8'd76, 1'b1, 1'b0};
3208: data_out = {8'd101, 8'd76, 1'b1, 1'b0};
3209: data_out = {8'd102, 8'd76, 1'b1, 1'b0};
3210: data_out = {8'd103, 8'd76, 1'b1, 1'b0};
3211: data_out = {8'd106, 8'd76, 1'b1, 1'b0};
3212: data_out = {8'd107, 8'd76, 1'b1, 1'b0};
3213: data_out = {8'd108, 8'd76, 1'b1, 1'b0};
3214: data_out = {8'd109, 8'd76, 1'b1, 1'b0};
3215: data_out = {8'd110, 8'd76, 1'b1, 1'b0};
3216: data_out = {8'd112, 8'd76, 1'b1, 1'b0};
3217: data_out = {8'd113, 8'd76, 1'b1, 1'b0};
3218: data_out = {8'd114, 8'd76, 1'b1, 1'b0};
3219: data_out = {8'd115, 8'd76, 1'b1, 1'b0};
3220: data_out = {8'd116, 8'd76, 1'b1, 1'b0};
3221: data_out = {8'd117, 8'd76, 1'b1, 1'b0};
3222: data_out = {8'd118, 8'd76, 1'b1, 1'b0};
3223: data_out = {8'd121, 8'd76, 1'b1, 1'b0};
3224: data_out = {8'd122, 8'd76, 1'b1, 1'b0};
3225: data_out = {8'd123, 8'd76, 1'b1, 1'b0};
3226: data_out = {8'd124, 8'd76, 1'b1, 1'b0};
3227: data_out = {8'd125, 8'd76, 1'b1, 1'b0};
3228: data_out = {8'd134, 8'd76, 1'b1, 1'b0};
3229: data_out = {8'd135, 8'd76, 1'b1, 1'b0};
3230: data_out = {8'd136, 8'd76, 1'b1, 1'b0};
3231: data_out = {8'd137, 8'd76, 1'b1, 1'b0};
3232: data_out = {8'd138, 8'd76, 1'b1, 1'b0};
3233: data_out = {8'd141, 8'd76, 1'b1, 1'b0};
3234: data_out = {8'd142, 8'd76, 1'b1, 1'b0};
3235: data_out = {8'd143, 8'd76, 1'b1, 1'b0};
3236: data_out = {8'd144, 8'd76, 1'b1, 1'b0};
3237: data_out = {8'd145, 8'd76, 1'b1, 1'b0};
3238: data_out = {8'd148, 8'd76, 1'b1, 1'b0};
3239: data_out = {8'd149, 8'd76, 1'b1, 1'b0};
3240: data_out = {8'd150, 8'd76, 1'b1, 1'b0};
3241: data_out = {8'd151, 8'd76, 1'b1, 1'b0};
3242: data_out = {8'd152, 8'd76, 1'b1, 1'b0};
3243: data_out = {8'd155, 8'd76, 1'b1, 1'b0};
3244: data_out = {8'd156, 8'd76, 1'b1, 1'b0};
3245: data_out = {8'd157, 8'd76, 1'b1, 1'b0};
3246: data_out = {8'd161, 8'd76, 1'b1, 1'b0};
3247: data_out = {8'd162, 8'd76, 1'b1, 1'b0};
3248: data_out = {8'd163, 8'd76, 1'b1, 1'b0};
3249: data_out = {8'd164, 8'd76, 1'b1, 1'b0};
3250: data_out = {8'd165, 8'd76, 1'b1, 1'b0};
3251: data_out = {8'd168, 8'd76, 1'b1, 1'b0};
3252: data_out = {8'd169, 8'd76, 1'b1, 1'b0};
3253: data_out = {8'd170, 8'd76, 1'b1, 1'b0};
3254: data_out = {8'd171, 8'd76, 1'b1, 1'b0};
3255: data_out = {8'd172, 8'd76, 1'b1, 1'b0};
3256: data_out = {8'd175, 8'd76, 1'b1, 1'b0};
3257: data_out = {8'd176, 8'd76, 1'b1, 1'b0};
3258: data_out = {8'd177, 8'd76, 1'b1, 1'b0};
3259: data_out = {8'd178, 8'd76, 1'b1, 1'b0};
3260: data_out = {8'd179, 8'd76, 1'b1, 1'b0};
3261: data_out = {8'd183, 8'd76, 1'b1, 1'b0};
3262: data_out = {8'd184, 8'd76, 1'b1, 1'b0};
3263: data_out = {8'd185, 8'd76, 1'b1, 1'b0};
3264: data_out = {8'd6, 8'd77, 1'b1, 1'b0};
3265: data_out = {8'd10, 8'd77, 1'b1, 1'b0};
3266: data_out = {8'd13, 8'd77, 1'b1, 1'b0};
3267: data_out = {8'd17, 8'd77, 1'b1, 1'b0};
3268: data_out = {8'd26, 8'd77, 1'b1, 1'b0};
3269: data_out = {8'd30, 8'd77, 1'b1, 1'b0};
3270: data_out = {8'd39, 8'd77, 1'b1, 1'b0};
3271: data_out = {8'd43, 8'd77, 1'b1, 1'b0};
3272: data_out = {8'd46, 8'd77, 1'b1, 1'b0};
3273: data_out = {8'd50, 8'd77, 1'b1, 1'b0};
3274: data_out = {8'd54, 8'd77, 1'b1, 1'b0};
3275: data_out = {8'd56, 8'd77, 1'b1, 1'b0};
3276: data_out = {8'd59, 8'd77, 1'b1, 1'b0};
3277: data_out = {8'd63, 8'd77, 1'b1, 1'b0};
3278: data_out = {8'd66, 8'd77, 1'b1, 1'b0};
3279: data_out = {8'd70, 8'd77, 1'b1, 1'b0};
3280: data_out = {8'd79, 8'd77, 1'b1, 1'b0};
3281: data_out = {8'd83, 8'd77, 1'b1, 1'b0};
3282: data_out = {8'd86, 8'd77, 1'b1, 1'b0};
3283: data_out = {8'd90, 8'd77, 1'b1, 1'b0};
3284: data_out = {8'd93, 8'd77, 1'b1, 1'b0};
3285: data_out = {8'd97, 8'd77, 1'b1, 1'b0};
3286: data_out = {8'd100, 8'd77, 1'b1, 1'b0};
3287: data_out = {8'd106, 8'd77, 1'b1, 1'b0};
3288: data_out = {8'd110, 8'd77, 1'b1, 1'b0};
3289: data_out = {8'd112, 8'd77, 1'b1, 1'b0};
3290: data_out = {8'd115, 8'd77, 1'b1, 1'b0};
3291: data_out = {8'd118, 8'd77, 1'b1, 1'b0};
3292: data_out = {8'd121, 8'd77, 1'b1, 1'b0};
3293: data_out = {8'd125, 8'd77, 1'b1, 1'b0};
3294: data_out = {8'd134, 8'd77, 1'b1, 1'b0};
3295: data_out = {8'd138, 8'd77, 1'b1, 1'b0};
3296: data_out = {8'd141, 8'd77, 1'b1, 1'b0};
3297: data_out = {8'd145, 8'd77, 1'b1, 1'b0};
3298: data_out = {8'd148, 8'd77, 1'b1, 1'b0};
3299: data_out = {8'd151, 8'd77, 1'b1, 1'b0};
3300: data_out = {8'd157, 8'd77, 1'b1, 1'b0};
3301: data_out = {8'd161, 8'd77, 1'b1, 1'b0};
3302: data_out = {8'd165, 8'd77, 1'b1, 1'b0};
3303: data_out = {8'd168, 8'd77, 1'b1, 1'b0};
3304: data_out = {8'd172, 8'd77, 1'b1, 1'b0};
3305: data_out = {8'd175, 8'd77, 1'b1, 1'b0};
3306: data_out = {8'd179, 8'd77, 1'b1, 1'b0};
3307: data_out = {8'd183, 8'd77, 1'b1, 1'b0};
3308: data_out = {8'd185, 8'd77, 1'b1, 1'b0};
3309: data_out = {8'd10, 8'd78, 1'b1, 1'b0};
3310: data_out = {8'd13, 8'd78, 1'b1, 1'b0};
3311: data_out = {8'd30, 8'd78, 1'b1, 1'b0};
3312: data_out = {8'd39, 8'd78, 1'b1, 1'b0};
3313: data_out = {8'd43, 8'd78, 1'b1, 1'b0};
3314: data_out = {8'd46, 8'd78, 1'b1, 1'b0};
3315: data_out = {8'd50, 8'd78, 1'b1, 1'b0};
3316: data_out = {8'd54, 8'd78, 1'b1, 1'b0};
3317: data_out = {8'd63, 8'd78, 1'b1, 1'b0};
3318: data_out = {8'd66, 8'd78, 1'b1, 1'b0};
3319: data_out = {8'd70, 8'd78, 1'b1, 1'b0};
3320: data_out = {8'd79, 8'd78, 1'b1, 1'b0};
3321: data_out = {8'd86, 8'd78, 1'b1, 1'b0};
3322: data_out = {8'd90, 8'd78, 1'b1, 1'b0};
3323: data_out = {8'd93, 8'd78, 1'b1, 1'b0};
3324: data_out = {8'd100, 8'd78, 1'b1, 1'b0};
3325: data_out = {8'd106, 8'd78, 1'b1, 1'b0};
3326: data_out = {8'd110, 8'd78, 1'b1, 1'b0};
3327: data_out = {8'd112, 8'd78, 1'b1, 1'b0};
3328: data_out = {8'd115, 8'd78, 1'b1, 1'b0};
3329: data_out = {8'd118, 8'd78, 1'b1, 1'b0};
3330: data_out = {8'd121, 8'd78, 1'b1, 1'b0};
3331: data_out = {8'd134, 8'd78, 1'b1, 1'b0};
3332: data_out = {8'd138, 8'd78, 1'b1, 1'b0};
3333: data_out = {8'd141, 8'd78, 1'b1, 1'b0};
3334: data_out = {8'd145, 8'd78, 1'b1, 1'b0};
3335: data_out = {8'd148, 8'd78, 1'b1, 1'b0};
3336: data_out = {8'd151, 8'd78, 1'b1, 1'b0};
3337: data_out = {8'd157, 8'd78, 1'b1, 1'b0};
3338: data_out = {8'd161, 8'd78, 1'b1, 1'b0};
3339: data_out = {8'd165, 8'd78, 1'b1, 1'b0};
3340: data_out = {8'd168, 8'd78, 1'b1, 1'b0};
3341: data_out = {8'd172, 8'd78, 1'b1, 1'b0};
3342: data_out = {8'd175, 8'd78, 1'b1, 1'b0};
3343: data_out = {8'd179, 8'd78, 1'b1, 1'b0};
3344: data_out = {8'd183, 8'd78, 1'b1, 1'b0};
3345: data_out = {8'd7, 8'd79, 1'b1, 1'b0};
3346: data_out = {8'd8, 8'd79, 1'b1, 1'b0};
3347: data_out = {8'd9, 8'd79, 1'b1, 1'b0};
3348: data_out = {8'd10, 8'd79, 1'b1, 1'b0};
3349: data_out = {8'd13, 8'd79, 1'b1, 1'b0};
3350: data_out = {8'd14, 8'd79, 1'b1, 1'b0};
3351: data_out = {8'd15, 8'd79, 1'b1, 1'b0};
3352: data_out = {8'd16, 8'd79, 1'b1, 1'b0};
3353: data_out = {8'd17, 8'd79, 1'b1, 1'b0};
3354: data_out = {8'd27, 8'd79, 1'b1, 1'b0};
3355: data_out = {8'd28, 8'd79, 1'b1, 1'b0};
3356: data_out = {8'd29, 8'd79, 1'b1, 1'b0};
3357: data_out = {8'd30, 8'd79, 1'b1, 1'b0};
3358: data_out = {8'd39, 8'd79, 1'b1, 1'b0};
3359: data_out = {8'd43, 8'd79, 1'b1, 1'b0};
3360: data_out = {8'd46, 8'd79, 1'b1, 1'b0};
3361: data_out = {8'd50, 8'd79, 1'b1, 1'b0};
3362: data_out = {8'd54, 8'd79, 1'b1, 1'b0};
3363: data_out = {8'd60, 8'd79, 1'b1, 1'b0};
3364: data_out = {8'd61, 8'd79, 1'b1, 1'b0};
3365: data_out = {8'd62, 8'd79, 1'b1, 1'b0};
3366: data_out = {8'd63, 8'd79, 1'b1, 1'b0};
3367: data_out = {8'd66, 8'd79, 1'b1, 1'b0};
3368: data_out = {8'd70, 8'd79, 1'b1, 1'b0};
3369: data_out = {8'd79, 8'd79, 1'b1, 1'b0};
3370: data_out = {8'd80, 8'd79, 1'b1, 1'b0};
3371: data_out = {8'd81, 8'd79, 1'b1, 1'b0};
3372: data_out = {8'd82, 8'd79, 1'b1, 1'b0};
3373: data_out = {8'd83, 8'd79, 1'b1, 1'b0};
3374: data_out = {8'd86, 8'd79, 1'b1, 1'b0};
3375: data_out = {8'd90, 8'd79, 1'b1, 1'b0};
3376: data_out = {8'd93, 8'd79, 1'b1, 1'b0};
3377: data_out = {8'd94, 8'd79, 1'b1, 1'b0};
3378: data_out = {8'd95, 8'd79, 1'b1, 1'b0};
3379: data_out = {8'd96, 8'd79, 1'b1, 1'b0};
3380: data_out = {8'd97, 8'd79, 1'b1, 1'b0};
3381: data_out = {8'd100, 8'd79, 1'b1, 1'b0};
3382: data_out = {8'd106, 8'd79, 1'b1, 1'b0};
3383: data_out = {8'd107, 8'd79, 1'b1, 1'b0};
3384: data_out = {8'd108, 8'd79, 1'b1, 1'b0};
3385: data_out = {8'd109, 8'd79, 1'b1, 1'b0};
3386: data_out = {8'd112, 8'd79, 1'b1, 1'b0};
3387: data_out = {8'd115, 8'd79, 1'b1, 1'b0};
3388: data_out = {8'd118, 8'd79, 1'b1, 1'b0};
3389: data_out = {8'd121, 8'd79, 1'b1, 1'b0};
3390: data_out = {8'd122, 8'd79, 1'b1, 1'b0};
3391: data_out = {8'd123, 8'd79, 1'b1, 1'b0};
3392: data_out = {8'd124, 8'd79, 1'b1, 1'b0};
3393: data_out = {8'd125, 8'd79, 1'b1, 1'b0};
3394: data_out = {8'd134, 8'd79, 1'b1, 1'b0};
3395: data_out = {8'd135, 8'd79, 1'b1, 1'b0};
3396: data_out = {8'd136, 8'd79, 1'b1, 1'b0};
3397: data_out = {8'd137, 8'd79, 1'b1, 1'b0};
3398: data_out = {8'd141, 8'd79, 1'b1, 1'b0};
3399: data_out = {8'd145, 8'd79, 1'b1, 1'b0};
3400: data_out = {8'd148, 8'd79, 1'b1, 1'b0};
3401: data_out = {8'd151, 8'd79, 1'b1, 1'b0};
3402: data_out = {8'd157, 8'd79, 1'b1, 1'b0};
3403: data_out = {8'd161, 8'd79, 1'b1, 1'b0};
3404: data_out = {8'd165, 8'd79, 1'b1, 1'b0};
3405: data_out = {8'd168, 8'd79, 1'b1, 1'b0};
3406: data_out = {8'd169, 8'd79, 1'b1, 1'b0};
3407: data_out = {8'd170, 8'd79, 1'b1, 1'b0};
3408: data_out = {8'd171, 8'd79, 1'b1, 1'b0};
3409: data_out = {8'd175, 8'd79, 1'b1, 1'b0};
3410: data_out = {8'd176, 8'd79, 1'b1, 1'b0};
3411: data_out = {8'd177, 8'd79, 1'b1, 1'b0};
3412: data_out = {8'd178, 8'd79, 1'b1, 1'b0};
3413: data_out = {8'd183, 8'd79, 1'b1, 1'b0};
3414: data_out = {8'd6, 8'd80, 1'b1, 1'b0};
3415: data_out = {8'd10, 8'd80, 1'b1, 1'b0};
3416: data_out = {8'd17, 8'd80, 1'b1, 1'b0};
3417: data_out = {8'd26, 8'd80, 1'b1, 1'b0};
3418: data_out = {8'd30, 8'd80, 1'b1, 1'b0};
3419: data_out = {8'd39, 8'd80, 1'b1, 1'b0};
3420: data_out = {8'd43, 8'd80, 1'b1, 1'b0};
3421: data_out = {8'd46, 8'd80, 1'b1, 1'b0};
3422: data_out = {8'd50, 8'd80, 1'b1, 1'b0};
3423: data_out = {8'd54, 8'd80, 1'b1, 1'b0};
3424: data_out = {8'd59, 8'd80, 1'b1, 1'b0};
3425: data_out = {8'd63, 8'd80, 1'b1, 1'b0};
3426: data_out = {8'd66, 8'd80, 1'b1, 1'b0};
3427: data_out = {8'd70, 8'd80, 1'b1, 1'b0};
3428: data_out = {8'd83, 8'd80, 1'b1, 1'b0};
3429: data_out = {8'd86, 8'd80, 1'b1, 1'b0};
3430: data_out = {8'd90, 8'd80, 1'b1, 1'b0};
3431: data_out = {8'd97, 8'd80, 1'b1, 1'b0};
3432: data_out = {8'd100, 8'd80, 1'b1, 1'b0};
3433: data_out = {8'd106, 8'd80, 1'b1, 1'b0};
3434: data_out = {8'd112, 8'd80, 1'b1, 1'b0};
3435: data_out = {8'd115, 8'd80, 1'b1, 1'b0};
3436: data_out = {8'd118, 8'd80, 1'b1, 1'b0};
3437: data_out = {8'd125, 8'd80, 1'b1, 1'b0};
3438: data_out = {8'd134, 8'd80, 1'b1, 1'b0};
3439: data_out = {8'd141, 8'd80, 1'b1, 1'b0};
3440: data_out = {8'd145, 8'd80, 1'b1, 1'b0};
3441: data_out = {8'd148, 8'd80, 1'b1, 1'b0};
3442: data_out = {8'd149, 8'd80, 1'b1, 1'b0};
3443: data_out = {8'd150, 8'd80, 1'b1, 1'b0};
3444: data_out = {8'd151, 8'd80, 1'b1, 1'b0};
3445: data_out = {8'd157, 8'd80, 1'b1, 1'b0};
3446: data_out = {8'd161, 8'd80, 1'b1, 1'b0};
3447: data_out = {8'd165, 8'd80, 1'b1, 1'b0};
3448: data_out = {8'd168, 8'd80, 1'b1, 1'b0};
3449: data_out = {8'd175, 8'd80, 1'b1, 1'b0};
3450: data_out = {8'd183, 8'd80, 1'b1, 1'b0};
3451: data_out = {8'd6, 8'd81, 1'b1, 1'b0};
3452: data_out = {8'd10, 8'd81, 1'b1, 1'b0};
3453: data_out = {8'd17, 8'd81, 1'b1, 1'b0};
3454: data_out = {8'd26, 8'd81, 1'b1, 1'b0};
3455: data_out = {8'd30, 8'd81, 1'b1, 1'b0};
3456: data_out = {8'd39, 8'd81, 1'b1, 1'b0};
3457: data_out = {8'd43, 8'd81, 1'b1, 1'b0};
3458: data_out = {8'd46, 8'd81, 1'b1, 1'b0};
3459: data_out = {8'd50, 8'd81, 1'b1, 1'b0};
3460: data_out = {8'd54, 8'd81, 1'b1, 1'b0};
3461: data_out = {8'd59, 8'd81, 1'b1, 1'b0};
3462: data_out = {8'd63, 8'd81, 1'b1, 1'b0};
3463: data_out = {8'd66, 8'd81, 1'b1, 1'b0};
3464: data_out = {8'd70, 8'd81, 1'b1, 1'b0};
3465: data_out = {8'd83, 8'd81, 1'b1, 1'b0};
3466: data_out = {8'd86, 8'd81, 1'b1, 1'b0};
3467: data_out = {8'd90, 8'd81, 1'b1, 1'b0};
3468: data_out = {8'd97, 8'd81, 1'b1, 1'b0};
3469: data_out = {8'd100, 8'd81, 1'b1, 1'b0};
3470: data_out = {8'd106, 8'd81, 1'b1, 1'b0};
3471: data_out = {8'd112, 8'd81, 1'b1, 1'b0};
3472: data_out = {8'd115, 8'd81, 1'b1, 1'b0};
3473: data_out = {8'd118, 8'd81, 1'b1, 1'b0};
3474: data_out = {8'd125, 8'd81, 1'b1, 1'b0};
3475: data_out = {8'd134, 8'd81, 1'b1, 1'b0};
3476: data_out = {8'd141, 8'd81, 1'b1, 1'b0};
3477: data_out = {8'd145, 8'd81, 1'b1, 1'b0};
3478: data_out = {8'd148, 8'd81, 1'b1, 1'b0};
3479: data_out = {8'd157, 8'd81, 1'b1, 1'b0};
3480: data_out = {8'd161, 8'd81, 1'b1, 1'b0};
3481: data_out = {8'd165, 8'd81, 1'b1, 1'b0};
3482: data_out = {8'd168, 8'd81, 1'b1, 1'b0};
3483: data_out = {8'd175, 8'd81, 1'b1, 1'b0};
3484: data_out = {8'd183, 8'd81, 1'b1, 1'b0};
3485: data_out = {8'd6, 8'd82, 1'b1, 1'b0};
3486: data_out = {8'd7, 8'd82, 1'b1, 1'b0};
3487: data_out = {8'd8, 8'd82, 1'b1, 1'b0};
3488: data_out = {8'd9, 8'd82, 1'b1, 1'b0};
3489: data_out = {8'd10, 8'd82, 1'b1, 1'b0};
3490: data_out = {8'd13, 8'd82, 1'b1, 1'b0};
3491: data_out = {8'd14, 8'd82, 1'b1, 1'b0};
3492: data_out = {8'd15, 8'd82, 1'b1, 1'b0};
3493: data_out = {8'd16, 8'd82, 1'b1, 1'b0};
3494: data_out = {8'd17, 8'd82, 1'b1, 1'b0};
3495: data_out = {8'd26, 8'd82, 1'b1, 1'b0};
3496: data_out = {8'd27, 8'd82, 1'b1, 1'b0};
3497: data_out = {8'd28, 8'd82, 1'b1, 1'b0};
3498: data_out = {8'd29, 8'd82, 1'b1, 1'b0};
3499: data_out = {8'd30, 8'd82, 1'b1, 1'b0};
3500: data_out = {8'd39, 8'd82, 1'b1, 1'b0};
3501: data_out = {8'd43, 8'd82, 1'b1, 1'b0};
3502: data_out = {8'd46, 8'd82, 1'b1, 1'b0};
3503: data_out = {8'd47, 8'd82, 1'b1, 1'b0};
3504: data_out = {8'd48, 8'd82, 1'b1, 1'b0};
3505: data_out = {8'd49, 8'd82, 1'b1, 1'b0};
3506: data_out = {8'd50, 8'd82, 1'b1, 1'b0};
3507: data_out = {8'd52, 8'd82, 1'b1, 1'b0};
3508: data_out = {8'd53, 8'd82, 1'b1, 1'b0};
3509: data_out = {8'd54, 8'd82, 1'b1, 1'b0};
3510: data_out = {8'd55, 8'd82, 1'b1, 1'b0};
3511: data_out = {8'd56, 8'd82, 1'b1, 1'b0};
3512: data_out = {8'd57, 8'd82, 1'b1, 1'b0};
3513: data_out = {8'd59, 8'd82, 1'b1, 1'b0};
3514: data_out = {8'd60, 8'd82, 1'b1, 1'b0};
3515: data_out = {8'd61, 8'd82, 1'b1, 1'b0};
3516: data_out = {8'd62, 8'd82, 1'b1, 1'b0};
3517: data_out = {8'd63, 8'd82, 1'b1, 1'b0};
3518: data_out = {8'd66, 8'd82, 1'b1, 1'b0};
3519: data_out = {8'd67, 8'd82, 1'b1, 1'b0};
3520: data_out = {8'd68, 8'd82, 1'b1, 1'b0};
3521: data_out = {8'd69, 8'd82, 1'b1, 1'b0};
3522: data_out = {8'd70, 8'd82, 1'b1, 1'b0};
3523: data_out = {8'd79, 8'd82, 1'b1, 1'b0};
3524: data_out = {8'd80, 8'd82, 1'b1, 1'b0};
3525: data_out = {8'd81, 8'd82, 1'b1, 1'b0};
3526: data_out = {8'd82, 8'd82, 1'b1, 1'b0};
3527: data_out = {8'd83, 8'd82, 1'b1, 1'b0};
3528: data_out = {8'd86, 8'd82, 1'b1, 1'b0};
3529: data_out = {8'd87, 8'd82, 1'b1, 1'b0};
3530: data_out = {8'd88, 8'd82, 1'b1, 1'b0};
3531: data_out = {8'd89, 8'd82, 1'b1, 1'b0};
3532: data_out = {8'd90, 8'd82, 1'b1, 1'b0};
3533: data_out = {8'd93, 8'd82, 1'b1, 1'b0};
3534: data_out = {8'd94, 8'd82, 1'b1, 1'b0};
3535: data_out = {8'd95, 8'd82, 1'b1, 1'b0};
3536: data_out = {8'd96, 8'd82, 1'b1, 1'b0};
3537: data_out = {8'd97, 8'd82, 1'b1, 1'b0};
3538: data_out = {8'd100, 8'd82, 1'b1, 1'b0};
3539: data_out = {8'd101, 8'd82, 1'b1, 1'b0};
3540: data_out = {8'd102, 8'd82, 1'b1, 1'b0};
3541: data_out = {8'd103, 8'd82, 1'b1, 1'b0};
3542: data_out = {8'd104, 8'd82, 1'b1, 1'b0};
3543: data_out = {8'd106, 8'd82, 1'b1, 1'b0};
3544: data_out = {8'd107, 8'd82, 1'b1, 1'b0};
3545: data_out = {8'd108, 8'd82, 1'b1, 1'b0};
3546: data_out = {8'd109, 8'd82, 1'b1, 1'b0};
3547: data_out = {8'd110, 8'd82, 1'b1, 1'b0};
3548: data_out = {8'd112, 8'd82, 1'b1, 1'b0};
3549: data_out = {8'd115, 8'd82, 1'b1, 1'b0};
3550: data_out = {8'd118, 8'd82, 1'b1, 1'b0};
3551: data_out = {8'd121, 8'd82, 1'b1, 1'b0};
3552: data_out = {8'd122, 8'd82, 1'b1, 1'b0};
3553: data_out = {8'd123, 8'd82, 1'b1, 1'b0};
3554: data_out = {8'd124, 8'd82, 1'b1, 1'b0};
3555: data_out = {8'd125, 8'd82, 1'b1, 1'b0};
3556: data_out = {8'd134, 8'd82, 1'b1, 1'b0};
3557: data_out = {8'd135, 8'd82, 1'b1, 1'b0};
3558: data_out = {8'd136, 8'd82, 1'b1, 1'b0};
3559: data_out = {8'd137, 8'd82, 1'b1, 1'b0};
3560: data_out = {8'd138, 8'd82, 1'b1, 1'b0};
3561: data_out = {8'd141, 8'd82, 1'b1, 1'b0};
3562: data_out = {8'd145, 8'd82, 1'b1, 1'b0};
3563: data_out = {8'd148, 8'd82, 1'b1, 1'b0};
3564: data_out = {8'd149, 8'd82, 1'b1, 1'b0};
3565: data_out = {8'd150, 8'd82, 1'b1, 1'b0};
3566: data_out = {8'd151, 8'd82, 1'b1, 1'b0};
3567: data_out = {8'd152, 8'd82, 1'b1, 1'b0};
3568: data_out = {8'd155, 8'd82, 1'b1, 1'b0};
3569: data_out = {8'd156, 8'd82, 1'b1, 1'b0};
3570: data_out = {8'd157, 8'd82, 1'b1, 1'b0};
3571: data_out = {8'd158, 8'd82, 1'b1, 1'b0};
3572: data_out = {8'd159, 8'd82, 1'b1, 1'b0};
3573: data_out = {8'd161, 8'd82, 1'b1, 1'b0};
3574: data_out = {8'd165, 8'd82, 1'b1, 1'b0};
3575: data_out = {8'd168, 8'd82, 1'b1, 1'b0};
3576: data_out = {8'd169, 8'd82, 1'b1, 1'b0};
3577: data_out = {8'd170, 8'd82, 1'b1, 1'b0};
3578: data_out = {8'd171, 8'd82, 1'b1, 1'b0};
3579: data_out = {8'd172, 8'd82, 1'b1, 1'b0};
3580: data_out = {8'd175, 8'd82, 1'b1, 1'b0};
3581: data_out = {8'd176, 8'd82, 1'b1, 1'b0};
3582: data_out = {8'd177, 8'd82, 1'b1, 1'b0};
3583: data_out = {8'd178, 8'd82, 1'b1, 1'b0};
3584: data_out = {8'd179, 8'd82, 1'b1, 1'b0};
3585: data_out = {8'd181, 8'd82, 1'b1, 1'b0};
3586: data_out = {8'd182, 8'd82, 1'b1, 1'b0};
3587: data_out = {8'd183, 8'd82, 1'b1, 1'b0};
3588: data_out = {8'd184, 8'd82, 1'b1, 1'b0};
3589: data_out = {8'd185, 8'd82, 1'b1, 1'b0};
3590: data_out = {8'd186, 8'd82, 1'b1, 1'b0};
3591: data_out = {8'd190, 8'd82, 1'b1, 1'b0};
3592: data_out = {8'd90, 8'd83, 1'b1, 1'b0};
3593: data_out = {8'd148, 8'd83, 1'b1, 1'b0};
3594: data_out = {8'd152, 8'd83, 1'b1, 1'b0};
3595: data_out = {8'd189, 8'd83, 1'b1, 1'b0};
3596: data_out = {8'd190, 8'd83, 1'b1, 1'b0};
3597: data_out = {8'd90, 8'd84, 1'b1, 1'b0};
3598: data_out = {8'd148, 8'd84, 1'b1, 1'b0};
3599: data_out = {8'd152, 8'd84, 1'b1, 1'b0};
3600: data_out = {8'd86, 8'd85, 1'b1, 1'b0};
3601: data_out = {8'd87, 8'd85, 1'b1, 1'b0};
3602: data_out = {8'd88, 8'd85, 1'b1, 1'b0};
3603: data_out = {8'd89, 8'd85, 1'b1, 1'b0};
3604: data_out = {8'd90, 8'd85, 1'b1, 1'b0};
3605: data_out = {8'd148, 8'd85, 1'b1, 1'b0};
3606: data_out = {8'd149, 8'd85, 1'b1, 1'b0};
3607: data_out = {8'd150, 8'd85, 1'b1, 1'b0};
3608: data_out = {8'd151, 8'd85, 1'b1, 1'b0};
3609: data_out = {8'd152, 8'd85, 1'b1, 1'b0};
3610: data_out = {8'd146, 8'd86, 1'b1, 1'b0};
3611: data_out = {8'd147, 8'd86, 1'b1, 1'b0};
3612: data_out = {8'd148, 8'd86, 1'b1, 1'b0};
3613: data_out = {8'd149, 8'd86, 1'b1, 1'b0};
3614: data_out = {8'd49, 8'd87, 1'b1, 1'b0};
3615: data_out = {8'd69, 8'd87, 1'b1, 1'b0};
3616: data_out = {8'd95, 8'd87, 1'b1, 1'b0};
3617: data_out = {8'd135, 8'd87, 1'b1, 1'b0};
3618: data_out = {8'd146, 8'd87, 1'b1, 1'b0};
3619: data_out = {8'd149, 8'd87, 1'b1, 1'b0};
3620: data_out = {8'd170, 8'd87, 1'b1, 1'b0};
3621: data_out = {8'd112, 8'd88, 1'b1, 1'b0};
3622: data_out = {8'd135, 8'd88, 1'b1, 1'b0};
3623: data_out = {8'd146, 8'd88, 1'b1, 1'b0};
3624: data_out = {8'd170, 8'd88, 1'b1, 1'b0};
3625: data_out = {8'd6, 8'd89, 1'b1, 1'b0};
3626: data_out = {8'd10, 8'd89, 1'b1, 1'b0};
3627: data_out = {8'd13, 8'd89, 1'b1, 1'b0};
3628: data_out = {8'd14, 8'd89, 1'b1, 1'b0};
3629: data_out = {8'd15, 8'd89, 1'b1, 1'b0};
3630: data_out = {8'd16, 8'd89, 1'b1, 1'b0};
3631: data_out = {8'd17, 8'd89, 1'b1, 1'b0};
3632: data_out = {8'd20, 8'd89, 1'b1, 1'b0};
3633: data_out = {8'd24, 8'd89, 1'b1, 1'b0};
3634: data_out = {8'd28, 8'd89, 1'b1, 1'b0};
3635: data_out = {8'd29, 8'd89, 1'b1, 1'b0};
3636: data_out = {8'd30, 8'd89, 1'b1, 1'b0};
3637: data_out = {8'd38, 8'd89, 1'b1, 1'b0};
3638: data_out = {8'd39, 8'd89, 1'b1, 1'b0};
3639: data_out = {8'd40, 8'd89, 1'b1, 1'b0};
3640: data_out = {8'd41, 8'd89, 1'b1, 1'b0};
3641: data_out = {8'd42, 8'd89, 1'b1, 1'b0};
3642: data_out = {8'd43, 8'd89, 1'b1, 1'b0};
3643: data_out = {8'd44, 8'd89, 1'b1, 1'b0};
3644: data_out = {8'd47, 8'd89, 1'b1, 1'b0};
3645: data_out = {8'd48, 8'd89, 1'b1, 1'b0};
3646: data_out = {8'd49, 8'd89, 1'b1, 1'b0};
3647: data_out = {8'd53, 8'd89, 1'b1, 1'b0};
3648: data_out = {8'd54, 8'd89, 1'b1, 1'b0};
3649: data_out = {8'd55, 8'd89, 1'b1, 1'b0};
3650: data_out = {8'd56, 8'd89, 1'b1, 1'b0};
3651: data_out = {8'd57, 8'd89, 1'b1, 1'b0};
3652: data_out = {8'd60, 8'd89, 1'b1, 1'b0};
3653: data_out = {8'd61, 8'd89, 1'b1, 1'b0};
3654: data_out = {8'd62, 8'd89, 1'b1, 1'b0};
3655: data_out = {8'd63, 8'd89, 1'b1, 1'b0};
3656: data_out = {8'd64, 8'd89, 1'b1, 1'b0};
3657: data_out = {8'd67, 8'd89, 1'b1, 1'b0};
3658: data_out = {8'd68, 8'd89, 1'b1, 1'b0};
3659: data_out = {8'd69, 8'd89, 1'b1, 1'b0};
3660: data_out = {8'd73, 8'd89, 1'b1, 1'b0};
3661: data_out = {8'd74, 8'd89, 1'b1, 1'b0};
3662: data_out = {8'd75, 8'd89, 1'b1, 1'b0};
3663: data_out = {8'd76, 8'd89, 1'b1, 1'b0};
3664: data_out = {8'd77, 8'd89, 1'b1, 1'b0};
3665: data_out = {8'd80, 8'd89, 1'b1, 1'b0};
3666: data_out = {8'd81, 8'd89, 1'b1, 1'b0};
3667: data_out = {8'd82, 8'd89, 1'b1, 1'b0};
3668: data_out = {8'd83, 8'd89, 1'b1, 1'b0};
3669: data_out = {8'd84, 8'd89, 1'b1, 1'b0};
3670: data_out = {8'd93, 8'd89, 1'b1, 1'b0};
3671: data_out = {8'd94, 8'd89, 1'b1, 1'b0};
3672: data_out = {8'd95, 8'd89, 1'b1, 1'b0};
3673: data_out = {8'd99, 8'd89, 1'b1, 1'b0};
3674: data_out = {8'd100, 8'd89, 1'b1, 1'b0};
3675: data_out = {8'd101, 8'd89, 1'b1, 1'b0};
3676: data_out = {8'd102, 8'd89, 1'b1, 1'b0};
3677: data_out = {8'd103, 8'd89, 1'b1, 1'b0};
3678: data_out = {8'd111, 8'd89, 1'b1, 1'b0};
3679: data_out = {8'd112, 8'd89, 1'b1, 1'b0};
3680: data_out = {8'd113, 8'd89, 1'b1, 1'b0};
3681: data_out = {8'd114, 8'd89, 1'b1, 1'b0};
3682: data_out = {8'd115, 8'd89, 1'b1, 1'b0};
3683: data_out = {8'd118, 8'd89, 1'b1, 1'b0};
3684: data_out = {8'd119, 8'd89, 1'b1, 1'b0};
3685: data_out = {8'd120, 8'd89, 1'b1, 1'b0};
3686: data_out = {8'd121, 8'd89, 1'b1, 1'b0};
3687: data_out = {8'd122, 8'd89, 1'b1, 1'b0};
3688: data_out = {8'd131, 8'd89, 1'b1, 1'b0};
3689: data_out = {8'd132, 8'd89, 1'b1, 1'b0};
3690: data_out = {8'd133, 8'd89, 1'b1, 1'b0};
3691: data_out = {8'd134, 8'd89, 1'b1, 1'b0};
3692: data_out = {8'd135, 8'd89, 1'b1, 1'b0};
3693: data_out = {8'd138, 8'd89, 1'b1, 1'b0};
3694: data_out = {8'd139, 8'd89, 1'b1, 1'b0};
3695: data_out = {8'd140, 8'd89, 1'b1, 1'b0};
3696: data_out = {8'd141, 8'd89, 1'b1, 1'b0};
3697: data_out = {8'd142, 8'd89, 1'b1, 1'b0};
3698: data_out = {8'd144, 8'd89, 1'b1, 1'b0};
3699: data_out = {8'd145, 8'd89, 1'b1, 1'b0};
3700: data_out = {8'd146, 8'd89, 1'b1, 1'b0};
3701: data_out = {8'd147, 8'd89, 1'b1, 1'b0};
3702: data_out = {8'd148, 8'd89, 1'b1, 1'b0};
3703: data_out = {8'd149, 8'd89, 1'b1, 1'b0};
3704: data_out = {8'd152, 8'd89, 1'b1, 1'b0};
3705: data_out = {8'd153, 8'd89, 1'b1, 1'b0};
3706: data_out = {8'd154, 8'd89, 1'b1, 1'b0};
3707: data_out = {8'd155, 8'd89, 1'b1, 1'b0};
3708: data_out = {8'd156, 8'd89, 1'b1, 1'b0};
3709: data_out = {8'd159, 8'd89, 1'b1, 1'b0};
3710: data_out = {8'd160, 8'd89, 1'b1, 1'b0};
3711: data_out = {8'd161, 8'd89, 1'b1, 1'b0};
3712: data_out = {8'd162, 8'd89, 1'b1, 1'b0};
3713: data_out = {8'd163, 8'd89, 1'b1, 1'b0};
3714: data_out = {8'd166, 8'd89, 1'b1, 1'b0};
3715: data_out = {8'd167, 8'd89, 1'b1, 1'b0};
3716: data_out = {8'd168, 8'd89, 1'b1, 1'b0};
3717: data_out = {8'd169, 8'd89, 1'b1, 1'b0};
3718: data_out = {8'd170, 8'd89, 1'b1, 1'b0};
3719: data_out = {8'd6, 8'd90, 1'b1, 1'b0};
3720: data_out = {8'd10, 8'd90, 1'b1, 1'b0};
3721: data_out = {8'd13, 8'd90, 1'b1, 1'b0};
3722: data_out = {8'd17, 8'd90, 1'b1, 1'b0};
3723: data_out = {8'd20, 8'd90, 1'b1, 1'b0};
3724: data_out = {8'd24, 8'd90, 1'b1, 1'b0};
3725: data_out = {8'd28, 8'd90, 1'b1, 1'b0};
3726: data_out = {8'd30, 8'd90, 1'b1, 1'b0};
3727: data_out = {8'd38, 8'd90, 1'b1, 1'b0};
3728: data_out = {8'd41, 8'd90, 1'b1, 1'b0};
3729: data_out = {8'd44, 8'd90, 1'b1, 1'b0};
3730: data_out = {8'd49, 8'd90, 1'b1, 1'b0};
3731: data_out = {8'd53, 8'd90, 1'b1, 1'b0};
3732: data_out = {8'd57, 8'd90, 1'b1, 1'b0};
3733: data_out = {8'd60, 8'd90, 1'b1, 1'b0};
3734: data_out = {8'd64, 8'd90, 1'b1, 1'b0};
3735: data_out = {8'd69, 8'd90, 1'b1, 1'b0};
3736: data_out = {8'd73, 8'd90, 1'b1, 1'b0};
3737: data_out = {8'd77, 8'd90, 1'b1, 1'b0};
3738: data_out = {8'd80, 8'd90, 1'b1, 1'b0};
3739: data_out = {8'd84, 8'd90, 1'b1, 1'b0};
3740: data_out = {8'd95, 8'd90, 1'b1, 1'b0};
3741: data_out = {8'd99, 8'd90, 1'b1, 1'b0};
3742: data_out = {8'd103, 8'd90, 1'b1, 1'b0};
3743: data_out = {8'd112, 8'd90, 1'b1, 1'b0};
3744: data_out = {8'd118, 8'd90, 1'b1, 1'b0};
3745: data_out = {8'd122, 8'd90, 1'b1, 1'b0};
3746: data_out = {8'd131, 8'd90, 1'b1, 1'b0};
3747: data_out = {8'd135, 8'd90, 1'b1, 1'b0};
3748: data_out = {8'd138, 8'd90, 1'b1, 1'b0};
3749: data_out = {8'd142, 8'd90, 1'b1, 1'b0};
3750: data_out = {8'd146, 8'd90, 1'b1, 1'b0};
3751: data_out = {8'd152, 8'd90, 1'b1, 1'b0};
3752: data_out = {8'd156, 8'd90, 1'b1, 1'b0};
3753: data_out = {8'd159, 8'd90, 1'b1, 1'b0};
3754: data_out = {8'd163, 8'd90, 1'b1, 1'b0};
3755: data_out = {8'd166, 8'd90, 1'b1, 1'b0};
3756: data_out = {8'd170, 8'd90, 1'b1, 1'b0};
3757: data_out = {8'd6, 8'd91, 1'b1, 1'b0};
3758: data_out = {8'd10, 8'd91, 1'b1, 1'b0};
3759: data_out = {8'd13, 8'd91, 1'b1, 1'b0};
3760: data_out = {8'd17, 8'd91, 1'b1, 1'b0};
3761: data_out = {8'd20, 8'd91, 1'b1, 1'b0};
3762: data_out = {8'd24, 8'd91, 1'b1, 1'b0};
3763: data_out = {8'd28, 8'd91, 1'b1, 1'b0};
3764: data_out = {8'd38, 8'd91, 1'b1, 1'b0};
3765: data_out = {8'd41, 8'd91, 1'b1, 1'b0};
3766: data_out = {8'd44, 8'd91, 1'b1, 1'b0};
3767: data_out = {8'd49, 8'd91, 1'b1, 1'b0};
3768: data_out = {8'd53, 8'd91, 1'b1, 1'b0};
3769: data_out = {8'd60, 8'd91, 1'b1, 1'b0};
3770: data_out = {8'd69, 8'd91, 1'b1, 1'b0};
3771: data_out = {8'd73, 8'd91, 1'b1, 1'b0};
3772: data_out = {8'd77, 8'd91, 1'b1, 1'b0};
3773: data_out = {8'd80, 8'd91, 1'b1, 1'b0};
3774: data_out = {8'd84, 8'd91, 1'b1, 1'b0};
3775: data_out = {8'd95, 8'd91, 1'b1, 1'b0};
3776: data_out = {8'd99, 8'd91, 1'b1, 1'b0};
3777: data_out = {8'd112, 8'd91, 1'b1, 1'b0};
3778: data_out = {8'd118, 8'd91, 1'b1, 1'b0};
3779: data_out = {8'd122, 8'd91, 1'b1, 1'b0};
3780: data_out = {8'd131, 8'd91, 1'b1, 1'b0};
3781: data_out = {8'd135, 8'd91, 1'b1, 1'b0};
3782: data_out = {8'd138, 8'd91, 1'b1, 1'b0};
3783: data_out = {8'd142, 8'd91, 1'b1, 1'b0};
3784: data_out = {8'd146, 8'd91, 1'b1, 1'b0};
3785: data_out = {8'd152, 8'd91, 1'b1, 1'b0};
3786: data_out = {8'd156, 8'd91, 1'b1, 1'b0};
3787: data_out = {8'd159, 8'd91, 1'b1, 1'b0};
3788: data_out = {8'd163, 8'd91, 1'b1, 1'b0};
3789: data_out = {8'd166, 8'd91, 1'b1, 1'b0};
3790: data_out = {8'd170, 8'd91, 1'b1, 1'b0};
3791: data_out = {8'd6, 8'd92, 1'b1, 1'b0};
3792: data_out = {8'd10, 8'd92, 1'b1, 1'b0};
3793: data_out = {8'd13, 8'd92, 1'b1, 1'b0};
3794: data_out = {8'd17, 8'd92, 1'b1, 1'b0};
3795: data_out = {8'd20, 8'd92, 1'b1, 1'b0};
3796: data_out = {8'd24, 8'd92, 1'b1, 1'b0};
3797: data_out = {8'd28, 8'd92, 1'b1, 1'b0};
3798: data_out = {8'd38, 8'd92, 1'b1, 1'b0};
3799: data_out = {8'd41, 8'd92, 1'b1, 1'b0};
3800: data_out = {8'd44, 8'd92, 1'b1, 1'b0};
3801: data_out = {8'd49, 8'd92, 1'b1, 1'b0};
3802: data_out = {8'd53, 8'd92, 1'b1, 1'b0};
3803: data_out = {8'd54, 8'd92, 1'b1, 1'b0};
3804: data_out = {8'd55, 8'd92, 1'b1, 1'b0};
3805: data_out = {8'd56, 8'd92, 1'b1, 1'b0};
3806: data_out = {8'd57, 8'd92, 1'b1, 1'b0};
3807: data_out = {8'd60, 8'd92, 1'b1, 1'b0};
3808: data_out = {8'd61, 8'd92, 1'b1, 1'b0};
3809: data_out = {8'd62, 8'd92, 1'b1, 1'b0};
3810: data_out = {8'd63, 8'd92, 1'b1, 1'b0};
3811: data_out = {8'd64, 8'd92, 1'b1, 1'b0};
3812: data_out = {8'd69, 8'd92, 1'b1, 1'b0};
3813: data_out = {8'd73, 8'd92, 1'b1, 1'b0};
3814: data_out = {8'd77, 8'd92, 1'b1, 1'b0};
3815: data_out = {8'd80, 8'd92, 1'b1, 1'b0};
3816: data_out = {8'd84, 8'd92, 1'b1, 1'b0};
3817: data_out = {8'd95, 8'd92, 1'b1, 1'b0};
3818: data_out = {8'd99, 8'd92, 1'b1, 1'b0};
3819: data_out = {8'd100, 8'd92, 1'b1, 1'b0};
3820: data_out = {8'd101, 8'd92, 1'b1, 1'b0};
3821: data_out = {8'd102, 8'd92, 1'b1, 1'b0};
3822: data_out = {8'd103, 8'd92, 1'b1, 1'b0};
3823: data_out = {8'd112, 8'd92, 1'b1, 1'b0};
3824: data_out = {8'd118, 8'd92, 1'b1, 1'b0};
3825: data_out = {8'd122, 8'd92, 1'b1, 1'b0};
3826: data_out = {8'd131, 8'd92, 1'b1, 1'b0};
3827: data_out = {8'd135, 8'd92, 1'b1, 1'b0};
3828: data_out = {8'd138, 8'd92, 1'b1, 1'b0};
3829: data_out = {8'd139, 8'd92, 1'b1, 1'b0};
3830: data_out = {8'd140, 8'd92, 1'b1, 1'b0};
3831: data_out = {8'd141, 8'd92, 1'b1, 1'b0};
3832: data_out = {8'd146, 8'd92, 1'b1, 1'b0};
3833: data_out = {8'd152, 8'd92, 1'b1, 1'b0};
3834: data_out = {8'd153, 8'd92, 1'b1, 1'b0};
3835: data_out = {8'd154, 8'd92, 1'b1, 1'b0};
3836: data_out = {8'd155, 8'd92, 1'b1, 1'b0};
3837: data_out = {8'd159, 8'd92, 1'b1, 1'b0};
3838: data_out = {8'd163, 8'd92, 1'b1, 1'b0};
3839: data_out = {8'd166, 8'd92, 1'b1, 1'b0};
3840: data_out = {8'd170, 8'd92, 1'b1, 1'b0};
3841: data_out = {8'd6, 8'd93, 1'b1, 1'b0};
3842: data_out = {8'd10, 8'd93, 1'b1, 1'b0};
3843: data_out = {8'd13, 8'd93, 1'b1, 1'b0};
3844: data_out = {8'd17, 8'd93, 1'b1, 1'b0};
3845: data_out = {8'd20, 8'd93, 1'b1, 1'b0};
3846: data_out = {8'd24, 8'd93, 1'b1, 1'b0};
3847: data_out = {8'd28, 8'd93, 1'b1, 1'b0};
3848: data_out = {8'd38, 8'd93, 1'b1, 1'b0};
3849: data_out = {8'd41, 8'd93, 1'b1, 1'b0};
3850: data_out = {8'd44, 8'd93, 1'b1, 1'b0};
3851: data_out = {8'd49, 8'd93, 1'b1, 1'b0};
3852: data_out = {8'd57, 8'd93, 1'b1, 1'b0};
3853: data_out = {8'd64, 8'd93, 1'b1, 1'b0};
3854: data_out = {8'd69, 8'd93, 1'b1, 1'b0};
3855: data_out = {8'd73, 8'd93, 1'b1, 1'b0};
3856: data_out = {8'd77, 8'd93, 1'b1, 1'b0};
3857: data_out = {8'd80, 8'd93, 1'b1, 1'b0};
3858: data_out = {8'd84, 8'd93, 1'b1, 1'b0};
3859: data_out = {8'd95, 8'd93, 1'b1, 1'b0};
3860: data_out = {8'd103, 8'd93, 1'b1, 1'b0};
3861: data_out = {8'd112, 8'd93, 1'b1, 1'b0};
3862: data_out = {8'd118, 8'd93, 1'b1, 1'b0};
3863: data_out = {8'd122, 8'd93, 1'b1, 1'b0};
3864: data_out = {8'd131, 8'd93, 1'b1, 1'b0};
3865: data_out = {8'd135, 8'd93, 1'b1, 1'b0};
3866: data_out = {8'd138, 8'd93, 1'b1, 1'b0};
3867: data_out = {8'd146, 8'd93, 1'b1, 1'b0};
3868: data_out = {8'd152, 8'd93, 1'b1, 1'b0};
3869: data_out = {8'd159, 8'd93, 1'b1, 1'b0};
3870: data_out = {8'd163, 8'd93, 1'b1, 1'b0};
3871: data_out = {8'd166, 8'd93, 1'b1, 1'b0};
3872: data_out = {8'd170, 8'd93, 1'b1, 1'b0};
3873: data_out = {8'd6, 8'd94, 1'b1, 1'b0};
3874: data_out = {8'd10, 8'd94, 1'b1, 1'b0};
3875: data_out = {8'd13, 8'd94, 1'b1, 1'b0};
3876: data_out = {8'd17, 8'd94, 1'b1, 1'b0};
3877: data_out = {8'd20, 8'd94, 1'b1, 1'b0};
3878: data_out = {8'd24, 8'd94, 1'b1, 1'b0};
3879: data_out = {8'd28, 8'd94, 1'b1, 1'b0};
3880: data_out = {8'd38, 8'd94, 1'b1, 1'b0};
3881: data_out = {8'd41, 8'd94, 1'b1, 1'b0};
3882: data_out = {8'd44, 8'd94, 1'b1, 1'b0};
3883: data_out = {8'd49, 8'd94, 1'b1, 1'b0};
3884: data_out = {8'd57, 8'd94, 1'b1, 1'b0};
3885: data_out = {8'd64, 8'd94, 1'b1, 1'b0};
3886: data_out = {8'd69, 8'd94, 1'b1, 1'b0};
3887: data_out = {8'd73, 8'd94, 1'b1, 1'b0};
3888: data_out = {8'd77, 8'd94, 1'b1, 1'b0};
3889: data_out = {8'd80, 8'd94, 1'b1, 1'b0};
3890: data_out = {8'd84, 8'd94, 1'b1, 1'b0};
3891: data_out = {8'd95, 8'd94, 1'b1, 1'b0};
3892: data_out = {8'd103, 8'd94, 1'b1, 1'b0};
3893: data_out = {8'd112, 8'd94, 1'b1, 1'b0};
3894: data_out = {8'd118, 8'd94, 1'b1, 1'b0};
3895: data_out = {8'd122, 8'd94, 1'b1, 1'b0};
3896: data_out = {8'd131, 8'd94, 1'b1, 1'b0};
3897: data_out = {8'd135, 8'd94, 1'b1, 1'b0};
3898: data_out = {8'd138, 8'd94, 1'b1, 1'b0};
3899: data_out = {8'd146, 8'd94, 1'b1, 1'b0};
3900: data_out = {8'd152, 8'd94, 1'b1, 1'b0};
3901: data_out = {8'd159, 8'd94, 1'b1, 1'b0};
3902: data_out = {8'd163, 8'd94, 1'b1, 1'b0};
3903: data_out = {8'd166, 8'd94, 1'b1, 1'b0};
3904: data_out = {8'd170, 8'd94, 1'b1, 1'b0};
3905: data_out = {8'd6, 8'd95, 1'b1, 1'b0};
3906: data_out = {8'd7, 8'd95, 1'b1, 1'b0};
3907: data_out = {8'd8, 8'd95, 1'b1, 1'b0};
3908: data_out = {8'd9, 8'd95, 1'b1, 1'b0};
3909: data_out = {8'd10, 8'd95, 1'b1, 1'b0};
3910: data_out = {8'd13, 8'd95, 1'b1, 1'b0};
3911: data_out = {8'd14, 8'd95, 1'b1, 1'b0};
3912: data_out = {8'd15, 8'd95, 1'b1, 1'b0};
3913: data_out = {8'd16, 8'd95, 1'b1, 1'b0};
3914: data_out = {8'd17, 8'd95, 1'b1, 1'b0};
3915: data_out = {8'd20, 8'd95, 1'b1, 1'b0};
3916: data_out = {8'd21, 8'd95, 1'b1, 1'b0};
3917: data_out = {8'd22, 8'd95, 1'b1, 1'b0};
3918: data_out = {8'd23, 8'd95, 1'b1, 1'b0};
3919: data_out = {8'd24, 8'd95, 1'b1, 1'b0};
3920: data_out = {8'd26, 8'd95, 1'b1, 1'b0};
3921: data_out = {8'd27, 8'd95, 1'b1, 1'b0};
3922: data_out = {8'd28, 8'd95, 1'b1, 1'b0};
3923: data_out = {8'd29, 8'd95, 1'b1, 1'b0};
3924: data_out = {8'd30, 8'd95, 1'b1, 1'b0};
3925: data_out = {8'd31, 8'd95, 1'b1, 1'b0};
3926: data_out = {8'd38, 8'd95, 1'b1, 1'b0};
3927: data_out = {8'd41, 8'd95, 1'b1, 1'b0};
3928: data_out = {8'd44, 8'd95, 1'b1, 1'b0};
3929: data_out = {8'd47, 8'd95, 1'b1, 1'b0};
3930: data_out = {8'd48, 8'd95, 1'b1, 1'b0};
3931: data_out = {8'd49, 8'd95, 1'b1, 1'b0};
3932: data_out = {8'd50, 8'd95, 1'b1, 1'b0};
3933: data_out = {8'd51, 8'd95, 1'b1, 1'b0};
3934: data_out = {8'd53, 8'd95, 1'b1, 1'b0};
3935: data_out = {8'd54, 8'd95, 1'b1, 1'b0};
3936: data_out = {8'd55, 8'd95, 1'b1, 1'b0};
3937: data_out = {8'd56, 8'd95, 1'b1, 1'b0};
3938: data_out = {8'd57, 8'd95, 1'b1, 1'b0};
3939: data_out = {8'd60, 8'd95, 1'b1, 1'b0};
3940: data_out = {8'd61, 8'd95, 1'b1, 1'b0};
3941: data_out = {8'd62, 8'd95, 1'b1, 1'b0};
3942: data_out = {8'd63, 8'd95, 1'b1, 1'b0};
3943: data_out = {8'd64, 8'd95, 1'b1, 1'b0};
3944: data_out = {8'd67, 8'd95, 1'b1, 1'b0};
3945: data_out = {8'd68, 8'd95, 1'b1, 1'b0};
3946: data_out = {8'd69, 8'd95, 1'b1, 1'b0};
3947: data_out = {8'd70, 8'd95, 1'b1, 1'b0};
3948: data_out = {8'd71, 8'd95, 1'b1, 1'b0};
3949: data_out = {8'd73, 8'd95, 1'b1, 1'b0};
3950: data_out = {8'd74, 8'd95, 1'b1, 1'b0};
3951: data_out = {8'd75, 8'd95, 1'b1, 1'b0};
3952: data_out = {8'd76, 8'd95, 1'b1, 1'b0};
3953: data_out = {8'd77, 8'd95, 1'b1, 1'b0};
3954: data_out = {8'd80, 8'd95, 1'b1, 1'b0};
3955: data_out = {8'd84, 8'd95, 1'b1, 1'b0};
3956: data_out = {8'd93, 8'd95, 1'b1, 1'b0};
3957: data_out = {8'd94, 8'd95, 1'b1, 1'b0};
3958: data_out = {8'd95, 8'd95, 1'b1, 1'b0};
3959: data_out = {8'd96, 8'd95, 1'b1, 1'b0};
3960: data_out = {8'd97, 8'd95, 1'b1, 1'b0};
3961: data_out = {8'd99, 8'd95, 1'b1, 1'b0};
3962: data_out = {8'd100, 8'd95, 1'b1, 1'b0};
3963: data_out = {8'd101, 8'd95, 1'b1, 1'b0};
3964: data_out = {8'd102, 8'd95, 1'b1, 1'b0};
3965: data_out = {8'd103, 8'd95, 1'b1, 1'b0};
3966: data_out = {8'd112, 8'd95, 1'b1, 1'b0};
3967: data_out = {8'd113, 8'd95, 1'b1, 1'b0};
3968: data_out = {8'd114, 8'd95, 1'b1, 1'b0};
3969: data_out = {8'd115, 8'd95, 1'b1, 1'b0};
3970: data_out = {8'd116, 8'd95, 1'b1, 1'b0};
3971: data_out = {8'd118, 8'd95, 1'b1, 1'b0};
3972: data_out = {8'd119, 8'd95, 1'b1, 1'b0};
3973: data_out = {8'd120, 8'd95, 1'b1, 1'b0};
3974: data_out = {8'd121, 8'd95, 1'b1, 1'b0};
3975: data_out = {8'd122, 8'd95, 1'b1, 1'b0};
3976: data_out = {8'd131, 8'd95, 1'b1, 1'b0};
3977: data_out = {8'd132, 8'd95, 1'b1, 1'b0};
3978: data_out = {8'd133, 8'd95, 1'b1, 1'b0};
3979: data_out = {8'd134, 8'd95, 1'b1, 1'b0};
3980: data_out = {8'd135, 8'd95, 1'b1, 1'b0};
3981: data_out = {8'd138, 8'd95, 1'b1, 1'b0};
3982: data_out = {8'd139, 8'd95, 1'b1, 1'b0};
3983: data_out = {8'd140, 8'd95, 1'b1, 1'b0};
3984: data_out = {8'd141, 8'd95, 1'b1, 1'b0};
3985: data_out = {8'd142, 8'd95, 1'b1, 1'b0};
3986: data_out = {8'd144, 8'd95, 1'b1, 1'b0};
3987: data_out = {8'd145, 8'd95, 1'b1, 1'b0};
3988: data_out = {8'd146, 8'd95, 1'b1, 1'b0};
3989: data_out = {8'd147, 8'd95, 1'b1, 1'b0};
3990: data_out = {8'd148, 8'd95, 1'b1, 1'b0};
3991: data_out = {8'd149, 8'd95, 1'b1, 1'b0};
3992: data_out = {8'd152, 8'd95, 1'b1, 1'b0};
3993: data_out = {8'd153, 8'd95, 1'b1, 1'b0};
3994: data_out = {8'd154, 8'd95, 1'b1, 1'b0};
3995: data_out = {8'd155, 8'd95, 1'b1, 1'b0};
3996: data_out = {8'd156, 8'd95, 1'b1, 1'b0};
3997: data_out = {8'd159, 8'd95, 1'b1, 1'b0};
3998: data_out = {8'd163, 8'd95, 1'b1, 1'b0};
3999: data_out = {8'd166, 8'd95, 1'b1, 1'b0};
4000: data_out = {8'd167, 8'd95, 1'b1, 1'b0};
4001: data_out = {8'd168, 8'd95, 1'b1, 1'b0};
4002: data_out = {8'd169, 8'd95, 1'b1, 1'b0};
4003: data_out = {8'd170, 8'd95, 1'b1, 1'b0};
4004: data_out = {8'd10, 8'd96, 1'b1, 1'b0};
4005: data_out = {8'd10, 8'd97, 1'b1, 1'b0};
4006: data_out = {8'd6, 8'd98, 1'b1, 1'b0};
4007: data_out = {8'd7, 8'd98, 1'b1, 1'b0};
4008: data_out = {8'd8, 8'd98, 1'b1, 1'b0};
4009: data_out = {8'd9, 8'd98, 1'b1, 1'b0};
4010: data_out = {8'd10, 8'd98, 1'b1, 1'b0};
4011: data_out = {8'd125, 8'd99, 1'b1, 1'b0};
4012: data_out = {8'd126, 8'd99, 1'b1, 1'b0};
4013: data_out = {8'd127, 8'd99, 1'b1, 1'b0};
4014: data_out = {8'd128, 8'd99, 1'b1, 1'b0};
4015: data_out = {8'd12, 8'd100, 1'b1, 1'b0};
4016: data_out = {8'd48, 8'd100, 1'b1, 1'b0};
4017: data_out = {8'd69, 8'd100, 1'b1, 1'b0};
4018: data_out = {8'd125, 8'd100, 1'b1, 1'b0};
4019: data_out = {8'd128, 8'd100, 1'b1, 1'b0};
4020: data_out = {8'd6, 8'd101, 1'b1, 1'b0};
4021: data_out = {8'd12, 8'd101, 1'b1, 1'b0};
4022: data_out = {8'd52, 8'd101, 1'b1, 1'b0};
4023: data_out = {8'd69, 8'd101, 1'b1, 1'b0};
4024: data_out = {8'd85, 8'd101, 1'b1, 1'b0};
4025: data_out = {8'd98, 8'd101, 1'b1, 1'b0};
4026: data_out = {8'd125, 8'd101, 1'b1, 1'b0};
4027: data_out = {8'd5, 8'd102, 1'b1, 1'b0};
4028: data_out = {8'd6, 8'd102, 1'b1, 1'b0};
4029: data_out = {8'd7, 8'd102, 1'b1, 1'b0};
4030: data_out = {8'd8, 8'd102, 1'b1, 1'b0};
4031: data_out = {8'd9, 8'd102, 1'b1, 1'b0};
4032: data_out = {8'd12, 8'd102, 1'b1, 1'b0};
4033: data_out = {8'd13, 8'd102, 1'b1, 1'b0};
4034: data_out = {8'd14, 8'd102, 1'b1, 1'b0};
4035: data_out = {8'd15, 8'd102, 1'b1, 1'b0};
4036: data_out = {8'd16, 8'd102, 1'b1, 1'b0};
4037: data_out = {8'd19, 8'd102, 1'b1, 1'b0};
4038: data_out = {8'd20, 8'd102, 1'b1, 1'b0};
4039: data_out = {8'd21, 8'd102, 1'b1, 1'b0};
4040: data_out = {8'd22, 8'd102, 1'b1, 1'b0};
4041: data_out = {8'd23, 8'd102, 1'b1, 1'b0};
4042: data_out = {8'd32, 8'd102, 1'b1, 1'b0};
4043: data_out = {8'd36, 8'd102, 1'b1, 1'b0};
4044: data_out = {8'd39, 8'd102, 1'b1, 1'b0};
4045: data_out = {8'd40, 8'd102, 1'b1, 1'b0};
4046: data_out = {8'd41, 8'd102, 1'b1, 1'b0};
4047: data_out = {8'd42, 8'd102, 1'b1, 1'b0};
4048: data_out = {8'd43, 8'd102, 1'b1, 1'b0};
4049: data_out = {8'd46, 8'd102, 1'b1, 1'b0};
4050: data_out = {8'd47, 8'd102, 1'b1, 1'b0};
4051: data_out = {8'd48, 8'd102, 1'b1, 1'b0};
4052: data_out = {8'd51, 8'd102, 1'b1, 1'b0};
4053: data_out = {8'd52, 8'd102, 1'b1, 1'b0};
4054: data_out = {8'd53, 8'd102, 1'b1, 1'b0};
4055: data_out = {8'd54, 8'd102, 1'b1, 1'b0};
4056: data_out = {8'd55, 8'd102, 1'b1, 1'b0};
4057: data_out = {8'd58, 8'd102, 1'b1, 1'b0};
4058: data_out = {8'd59, 8'd102, 1'b1, 1'b0};
4059: data_out = {8'd60, 8'd102, 1'b1, 1'b0};
4060: data_out = {8'd61, 8'd102, 1'b1, 1'b0};
4061: data_out = {8'd62, 8'd102, 1'b1, 1'b0};
4062: data_out = {8'd65, 8'd102, 1'b1, 1'b0};
4063: data_out = {8'd66, 8'd102, 1'b1, 1'b0};
4064: data_out = {8'd67, 8'd102, 1'b1, 1'b0};
4065: data_out = {8'd68, 8'd102, 1'b1, 1'b0};
4066: data_out = {8'd69, 8'd102, 1'b1, 1'b0};
4067: data_out = {8'd78, 8'd102, 1'b1, 1'b0};
4068: data_out = {8'd79, 8'd102, 1'b1, 1'b0};
4069: data_out = {8'd80, 8'd102, 1'b1, 1'b0};
4070: data_out = {8'd81, 8'd102, 1'b1, 1'b0};
4071: data_out = {8'd82, 8'd102, 1'b1, 1'b0};
4072: data_out = {8'd84, 8'd102, 1'b1, 1'b0};
4073: data_out = {8'd85, 8'd102, 1'b1, 1'b0};
4074: data_out = {8'd86, 8'd102, 1'b1, 1'b0};
4075: data_out = {8'd87, 8'd102, 1'b1, 1'b0};
4076: data_out = {8'd88, 8'd102, 1'b1, 1'b0};
4077: data_out = {8'd91, 8'd102, 1'b1, 1'b0};
4078: data_out = {8'd92, 8'd102, 1'b1, 1'b0};
4079: data_out = {8'd93, 8'd102, 1'b1, 1'b0};
4080: data_out = {8'd94, 8'd102, 1'b1, 1'b0};
4081: data_out = {8'd95, 8'd102, 1'b1, 1'b0};
4082: data_out = {8'd97, 8'd102, 1'b1, 1'b0};
4083: data_out = {8'd98, 8'd102, 1'b1, 1'b0};
4084: data_out = {8'd99, 8'd102, 1'b1, 1'b0};
4085: data_out = {8'd100, 8'd102, 1'b1, 1'b0};
4086: data_out = {8'd101, 8'd102, 1'b1, 1'b0};
4087: data_out = {8'd104, 8'd102, 1'b1, 1'b0};
4088: data_out = {8'd105, 8'd102, 1'b1, 1'b0};
4089: data_out = {8'd106, 8'd102, 1'b1, 1'b0};
4090: data_out = {8'd107, 8'd102, 1'b1, 1'b0};
4091: data_out = {8'd108, 8'd102, 1'b1, 1'b0};
4092: data_out = {8'd111, 8'd102, 1'b1, 1'b0};
4093: data_out = {8'd112, 8'd102, 1'b1, 1'b0};
4094: data_out = {8'd113, 8'd102, 1'b1, 1'b0};
4095: data_out = {8'd114, 8'd102, 1'b1, 1'b0};
4096: data_out = {8'd115, 8'd102, 1'b1, 1'b0};
4097: data_out = {8'd123, 8'd102, 1'b1, 1'b0};
4098: data_out = {8'd124, 8'd102, 1'b1, 1'b0};
4099: data_out = {8'd125, 8'd102, 1'b1, 1'b0};
4100: data_out = {8'd126, 8'd102, 1'b1, 1'b0};
4101: data_out = {8'd127, 8'd102, 1'b1, 1'b0};
4102: data_out = {8'd128, 8'd102, 1'b1, 1'b0};
4103: data_out = {8'd132, 8'd102, 1'b1, 1'b0};
4104: data_out = {8'd133, 8'd102, 1'b1, 1'b0};
4105: data_out = {8'd134, 8'd102, 1'b1, 1'b0};
4106: data_out = {8'd137, 8'd102, 1'b1, 1'b0};
4107: data_out = {8'd138, 8'd102, 1'b1, 1'b0};
4108: data_out = {8'd139, 8'd102, 1'b1, 1'b0};
4109: data_out = {8'd140, 8'd102, 1'b1, 1'b0};
4110: data_out = {8'd141, 8'd102, 1'b1, 1'b0};
4111: data_out = {8'd143, 8'd102, 1'b1, 1'b0};
4112: data_out = {8'd144, 8'd102, 1'b1, 1'b0};
4113: data_out = {8'd145, 8'd102, 1'b1, 1'b0};
4114: data_out = {8'd146, 8'd102, 1'b1, 1'b0};
4115: data_out = {8'd147, 8'd102, 1'b1, 1'b0};
4116: data_out = {8'd148, 8'd102, 1'b1, 1'b0};
4117: data_out = {8'd149, 8'd102, 1'b1, 1'b0};
4118: data_out = {8'd6, 8'd103, 1'b1, 1'b0};
4119: data_out = {8'd12, 8'd103, 1'b1, 1'b0};
4120: data_out = {8'd16, 8'd103, 1'b1, 1'b0};
4121: data_out = {8'd19, 8'd103, 1'b1, 1'b0};
4122: data_out = {8'd23, 8'd103, 1'b1, 1'b0};
4123: data_out = {8'd32, 8'd103, 1'b1, 1'b0};
4124: data_out = {8'd36, 8'd103, 1'b1, 1'b0};
4125: data_out = {8'd39, 8'd103, 1'b1, 1'b0};
4126: data_out = {8'd43, 8'd103, 1'b1, 1'b0};
4127: data_out = {8'd48, 8'd103, 1'b1, 1'b0};
4128: data_out = {8'd52, 8'd103, 1'b1, 1'b0};
4129: data_out = {8'd58, 8'd103, 1'b1, 1'b0};
4130: data_out = {8'd62, 8'd103, 1'b1, 1'b0};
4131: data_out = {8'd65, 8'd103, 1'b1, 1'b0};
4132: data_out = {8'd69, 8'd103, 1'b1, 1'b0};
4133: data_out = {8'd78, 8'd103, 1'b1, 1'b0};
4134: data_out = {8'd82, 8'd103, 1'b1, 1'b0};
4135: data_out = {8'd85, 8'd103, 1'b1, 1'b0};
4136: data_out = {8'd91, 8'd103, 1'b1, 1'b0};
4137: data_out = {8'd95, 8'd103, 1'b1, 1'b0};
4138: data_out = {8'd98, 8'd103, 1'b1, 1'b0};
4139: data_out = {8'd104, 8'd103, 1'b1, 1'b0};
4140: data_out = {8'd108, 8'd103, 1'b1, 1'b0};
4141: data_out = {8'd111, 8'd103, 1'b1, 1'b0};
4142: data_out = {8'd115, 8'd103, 1'b1, 1'b0};
4143: data_out = {8'd125, 8'd103, 1'b1, 1'b0};
4144: data_out = {8'd132, 8'd103, 1'b1, 1'b0};
4145: data_out = {8'd134, 8'd103, 1'b1, 1'b0};
4146: data_out = {8'd137, 8'd103, 1'b1, 1'b0};
4147: data_out = {8'd141, 8'd103, 1'b1, 1'b0};
4148: data_out = {8'd143, 8'd103, 1'b1, 1'b0};
4149: data_out = {8'd146, 8'd103, 1'b1, 1'b0};
4150: data_out = {8'd149, 8'd103, 1'b1, 1'b0};
4151: data_out = {8'd6, 8'd104, 1'b1, 1'b0};
4152: data_out = {8'd12, 8'd104, 1'b1, 1'b0};
4153: data_out = {8'd16, 8'd104, 1'b1, 1'b0};
4154: data_out = {8'd19, 8'd104, 1'b1, 1'b0};
4155: data_out = {8'd23, 8'd104, 1'b1, 1'b0};
4156: data_out = {8'd32, 8'd104, 1'b1, 1'b0};
4157: data_out = {8'd36, 8'd104, 1'b1, 1'b0};
4158: data_out = {8'd39, 8'd104, 1'b1, 1'b0};
4159: data_out = {8'd43, 8'd104, 1'b1, 1'b0};
4160: data_out = {8'd48, 8'd104, 1'b1, 1'b0};
4161: data_out = {8'd52, 8'd104, 1'b1, 1'b0};
4162: data_out = {8'd58, 8'd104, 1'b1, 1'b0};
4163: data_out = {8'd62, 8'd104, 1'b1, 1'b0};
4164: data_out = {8'd65, 8'd104, 1'b1, 1'b0};
4165: data_out = {8'd69, 8'd104, 1'b1, 1'b0};
4166: data_out = {8'd78, 8'd104, 1'b1, 1'b0};
4167: data_out = {8'd85, 8'd104, 1'b1, 1'b0};
4168: data_out = {8'd95, 8'd104, 1'b1, 1'b0};
4169: data_out = {8'd98, 8'd104, 1'b1, 1'b0};
4170: data_out = {8'd104, 8'd104, 1'b1, 1'b0};
4171: data_out = {8'd108, 8'd104, 1'b1, 1'b0};
4172: data_out = {8'd111, 8'd104, 1'b1, 1'b0};
4173: data_out = {8'd125, 8'd104, 1'b1, 1'b0};
4174: data_out = {8'd132, 8'd104, 1'b1, 1'b0};
4175: data_out = {8'd137, 8'd104, 1'b1, 1'b0};
4176: data_out = {8'd141, 8'd104, 1'b1, 1'b0};
4177: data_out = {8'd143, 8'd104, 1'b1, 1'b0};
4178: data_out = {8'd146, 8'd104, 1'b1, 1'b0};
4179: data_out = {8'd149, 8'd104, 1'b1, 1'b0};
4180: data_out = {8'd6, 8'd105, 1'b1, 1'b0};
4181: data_out = {8'd12, 8'd105, 1'b1, 1'b0};
4182: data_out = {8'd16, 8'd105, 1'b1, 1'b0};
4183: data_out = {8'd19, 8'd105, 1'b1, 1'b0};
4184: data_out = {8'd20, 8'd105, 1'b1, 1'b0};
4185: data_out = {8'd21, 8'd105, 1'b1, 1'b0};
4186: data_out = {8'd22, 8'd105, 1'b1, 1'b0};
4187: data_out = {8'd32, 8'd105, 1'b1, 1'b0};
4188: data_out = {8'd36, 8'd105, 1'b1, 1'b0};
4189: data_out = {8'd39, 8'd105, 1'b1, 1'b0};
4190: data_out = {8'd43, 8'd105, 1'b1, 1'b0};
4191: data_out = {8'd48, 8'd105, 1'b1, 1'b0};
4192: data_out = {8'd52, 8'd105, 1'b1, 1'b0};
4193: data_out = {8'd58, 8'd105, 1'b1, 1'b0};
4194: data_out = {8'd59, 8'd105, 1'b1, 1'b0};
4195: data_out = {8'd60, 8'd105, 1'b1, 1'b0};
4196: data_out = {8'd61, 8'd105, 1'b1, 1'b0};
4197: data_out = {8'd65, 8'd105, 1'b1, 1'b0};
4198: data_out = {8'd69, 8'd105, 1'b1, 1'b0};
4199: data_out = {8'd78, 8'd105, 1'b1, 1'b0};
4200: data_out = {8'd79, 8'd105, 1'b1, 1'b0};
4201: data_out = {8'd80, 8'd105, 1'b1, 1'b0};
4202: data_out = {8'd81, 8'd105, 1'b1, 1'b0};
4203: data_out = {8'd82, 8'd105, 1'b1, 1'b0};
4204: data_out = {8'd85, 8'd105, 1'b1, 1'b0};
4205: data_out = {8'd92, 8'd105, 1'b1, 1'b0};
4206: data_out = {8'd93, 8'd105, 1'b1, 1'b0};
4207: data_out = {8'd94, 8'd105, 1'b1, 1'b0};
4208: data_out = {8'd95, 8'd105, 1'b1, 1'b0};
4209: data_out = {8'd98, 8'd105, 1'b1, 1'b0};
4210: data_out = {8'd104, 8'd105, 1'b1, 1'b0};
4211: data_out = {8'd105, 8'd105, 1'b1, 1'b0};
4212: data_out = {8'd106, 8'd105, 1'b1, 1'b0};
4213: data_out = {8'd107, 8'd105, 1'b1, 1'b0};
4214: data_out = {8'd111, 8'd105, 1'b1, 1'b0};
4215: data_out = {8'd112, 8'd105, 1'b1, 1'b0};
4216: data_out = {8'd113, 8'd105, 1'b1, 1'b0};
4217: data_out = {8'd114, 8'd105, 1'b1, 1'b0};
4218: data_out = {8'd115, 8'd105, 1'b1, 1'b0};
4219: data_out = {8'd125, 8'd105, 1'b1, 1'b0};
4220: data_out = {8'd132, 8'd105, 1'b1, 1'b0};
4221: data_out = {8'd137, 8'd105, 1'b1, 1'b0};
4222: data_out = {8'd141, 8'd105, 1'b1, 1'b0};
4223: data_out = {8'd143, 8'd105, 1'b1, 1'b0};
4224: data_out = {8'd146, 8'd105, 1'b1, 1'b0};
4225: data_out = {8'd149, 8'd105, 1'b1, 1'b0};
4226: data_out = {8'd6, 8'd106, 1'b1, 1'b0};
4227: data_out = {8'd12, 8'd106, 1'b1, 1'b0};
4228: data_out = {8'd16, 8'd106, 1'b1, 1'b0};
4229: data_out = {8'd19, 8'd106, 1'b1, 1'b0};
4230: data_out = {8'd32, 8'd106, 1'b1, 1'b0};
4231: data_out = {8'd36, 8'd106, 1'b1, 1'b0};
4232: data_out = {8'd39, 8'd106, 1'b1, 1'b0};
4233: data_out = {8'd43, 8'd106, 1'b1, 1'b0};
4234: data_out = {8'd48, 8'd106, 1'b1, 1'b0};
4235: data_out = {8'd52, 8'd106, 1'b1, 1'b0};
4236: data_out = {8'd58, 8'd106, 1'b1, 1'b0};
4237: data_out = {8'd65, 8'd106, 1'b1, 1'b0};
4238: data_out = {8'd69, 8'd106, 1'b1, 1'b0};
4239: data_out = {8'd82, 8'd106, 1'b1, 1'b0};
4240: data_out = {8'd85, 8'd106, 1'b1, 1'b0};
4241: data_out = {8'd91, 8'd106, 1'b1, 1'b0};
4242: data_out = {8'd95, 8'd106, 1'b1, 1'b0};
4243: data_out = {8'd98, 8'd106, 1'b1, 1'b0};
4244: data_out = {8'd104, 8'd106, 1'b1, 1'b0};
4245: data_out = {8'd115, 8'd106, 1'b1, 1'b0};
4246: data_out = {8'd125, 8'd106, 1'b1, 1'b0};
4247: data_out = {8'd132, 8'd106, 1'b1, 1'b0};
4248: data_out = {8'd137, 8'd106, 1'b1, 1'b0};
4249: data_out = {8'd141, 8'd106, 1'b1, 1'b0};
4250: data_out = {8'd143, 8'd106, 1'b1, 1'b0};
4251: data_out = {8'd146, 8'd106, 1'b1, 1'b0};
4252: data_out = {8'd149, 8'd106, 1'b1, 1'b0};
4253: data_out = {8'd6, 8'd107, 1'b1, 1'b0};
4254: data_out = {8'd12, 8'd107, 1'b1, 1'b0};
4255: data_out = {8'd16, 8'd107, 1'b1, 1'b0};
4256: data_out = {8'd19, 8'd107, 1'b1, 1'b0};
4257: data_out = {8'd32, 8'd107, 1'b1, 1'b0};
4258: data_out = {8'd36, 8'd107, 1'b1, 1'b0};
4259: data_out = {8'd39, 8'd107, 1'b1, 1'b0};
4260: data_out = {8'd43, 8'd107, 1'b1, 1'b0};
4261: data_out = {8'd48, 8'd107, 1'b1, 1'b0};
4262: data_out = {8'd52, 8'd107, 1'b1, 1'b0};
4263: data_out = {8'd58, 8'd107, 1'b1, 1'b0};
4264: data_out = {8'd65, 8'd107, 1'b1, 1'b0};
4265: data_out = {8'd69, 8'd107, 1'b1, 1'b0};
4266: data_out = {8'd82, 8'd107, 1'b1, 1'b0};
4267: data_out = {8'd85, 8'd107, 1'b1, 1'b0};
4268: data_out = {8'd91, 8'd107, 1'b1, 1'b0};
4269: data_out = {8'd95, 8'd107, 1'b1, 1'b0};
4270: data_out = {8'd98, 8'd107, 1'b1, 1'b0};
4271: data_out = {8'd104, 8'd107, 1'b1, 1'b0};
4272: data_out = {8'd115, 8'd107, 1'b1, 1'b0};
4273: data_out = {8'd125, 8'd107, 1'b1, 1'b0};
4274: data_out = {8'd132, 8'd107, 1'b1, 1'b0};
4275: data_out = {8'd137, 8'd107, 1'b1, 1'b0};
4276: data_out = {8'd141, 8'd107, 1'b1, 1'b0};
4277: data_out = {8'd143, 8'd107, 1'b1, 1'b0};
4278: data_out = {8'd146, 8'd107, 1'b1, 1'b0};
4279: data_out = {8'd149, 8'd107, 1'b1, 1'b0};
4280: data_out = {8'd6, 8'd108, 1'b1, 1'b0};
4281: data_out = {8'd7, 8'd108, 1'b1, 1'b0};
4282: data_out = {8'd8, 8'd108, 1'b1, 1'b0};
4283: data_out = {8'd9, 8'd108, 1'b1, 1'b0};
4284: data_out = {8'd10, 8'd108, 1'b1, 1'b0};
4285: data_out = {8'd12, 8'd108, 1'b1, 1'b0};
4286: data_out = {8'd16, 8'd108, 1'b1, 1'b0};
4287: data_out = {8'd19, 8'd108, 1'b1, 1'b0};
4288: data_out = {8'd20, 8'd108, 1'b1, 1'b0};
4289: data_out = {8'd21, 8'd108, 1'b1, 1'b0};
4290: data_out = {8'd22, 8'd108, 1'b1, 1'b0};
4291: data_out = {8'd23, 8'd108, 1'b1, 1'b0};
4292: data_out = {8'd32, 8'd108, 1'b1, 1'b0};
4293: data_out = {8'd33, 8'd108, 1'b1, 1'b0};
4294: data_out = {8'd34, 8'd108, 1'b1, 1'b0};
4295: data_out = {8'd35, 8'd108, 1'b1, 1'b0};
4296: data_out = {8'd36, 8'd108, 1'b1, 1'b0};
4297: data_out = {8'd39, 8'd108, 1'b1, 1'b0};
4298: data_out = {8'd43, 8'd108, 1'b1, 1'b0};
4299: data_out = {8'd46, 8'd108, 1'b1, 1'b0};
4300: data_out = {8'd47, 8'd108, 1'b1, 1'b0};
4301: data_out = {8'd48, 8'd108, 1'b1, 1'b0};
4302: data_out = {8'd49, 8'd108, 1'b1, 1'b0};
4303: data_out = {8'd50, 8'd108, 1'b1, 1'b0};
4304: data_out = {8'd52, 8'd108, 1'b1, 1'b0};
4305: data_out = {8'd53, 8'd108, 1'b1, 1'b0};
4306: data_out = {8'd54, 8'd108, 1'b1, 1'b0};
4307: data_out = {8'd55, 8'd108, 1'b1, 1'b0};
4308: data_out = {8'd56, 8'd108, 1'b1, 1'b0};
4309: data_out = {8'd58, 8'd108, 1'b1, 1'b0};
4310: data_out = {8'd59, 8'd108, 1'b1, 1'b0};
4311: data_out = {8'd60, 8'd108, 1'b1, 1'b0};
4312: data_out = {8'd61, 8'd108, 1'b1, 1'b0};
4313: data_out = {8'd62, 8'd108, 1'b1, 1'b0};
4314: data_out = {8'd65, 8'd108, 1'b1, 1'b0};
4315: data_out = {8'd66, 8'd108, 1'b1, 1'b0};
4316: data_out = {8'd67, 8'd108, 1'b1, 1'b0};
4317: data_out = {8'd68, 8'd108, 1'b1, 1'b0};
4318: data_out = {8'd69, 8'd108, 1'b1, 1'b0};
4319: data_out = {8'd78, 8'd108, 1'b1, 1'b0};
4320: data_out = {8'd79, 8'd108, 1'b1, 1'b0};
4321: data_out = {8'd80, 8'd108, 1'b1, 1'b0};
4322: data_out = {8'd81, 8'd108, 1'b1, 1'b0};
4323: data_out = {8'd82, 8'd108, 1'b1, 1'b0};
4324: data_out = {8'd85, 8'd108, 1'b1, 1'b0};
4325: data_out = {8'd86, 8'd108, 1'b1, 1'b0};
4326: data_out = {8'd87, 8'd108, 1'b1, 1'b0};
4327: data_out = {8'd88, 8'd108, 1'b1, 1'b0};
4328: data_out = {8'd89, 8'd108, 1'b1, 1'b0};
4329: data_out = {8'd91, 8'd108, 1'b1, 1'b0};
4330: data_out = {8'd92, 8'd108, 1'b1, 1'b0};
4331: data_out = {8'd93, 8'd108, 1'b1, 1'b0};
4332: data_out = {8'd94, 8'd108, 1'b1, 1'b0};
4333: data_out = {8'd95, 8'd108, 1'b1, 1'b0};
4334: data_out = {8'd98, 8'd108, 1'b1, 1'b0};
4335: data_out = {8'd99, 8'd108, 1'b1, 1'b0};
4336: data_out = {8'd100, 8'd108, 1'b1, 1'b0};
4337: data_out = {8'd101, 8'd108, 1'b1, 1'b0};
4338: data_out = {8'd102, 8'd108, 1'b1, 1'b0};
4339: data_out = {8'd104, 8'd108, 1'b1, 1'b0};
4340: data_out = {8'd105, 8'd108, 1'b1, 1'b0};
4341: data_out = {8'd106, 8'd108, 1'b1, 1'b0};
4342: data_out = {8'd107, 8'd108, 1'b1, 1'b0};
4343: data_out = {8'd108, 8'd108, 1'b1, 1'b0};
4344: data_out = {8'd111, 8'd108, 1'b1, 1'b0};
4345: data_out = {8'd112, 8'd108, 1'b1, 1'b0};
4346: data_out = {8'd113, 8'd108, 1'b1, 1'b0};
4347: data_out = {8'd114, 8'd108, 1'b1, 1'b0};
4348: data_out = {8'd115, 8'd108, 1'b1, 1'b0};
4349: data_out = {8'd123, 8'd108, 1'b1, 1'b0};
4350: data_out = {8'd124, 8'd108, 1'b1, 1'b0};
4351: data_out = {8'd125, 8'd108, 1'b1, 1'b0};
4352: data_out = {8'd126, 8'd108, 1'b1, 1'b0};
4353: data_out = {8'd127, 8'd108, 1'b1, 1'b0};
4354: data_out = {8'd128, 8'd108, 1'b1, 1'b0};
4355: data_out = {8'd130, 8'd108, 1'b1, 1'b0};
4356: data_out = {8'd131, 8'd108, 1'b1, 1'b0};
4357: data_out = {8'd132, 8'd108, 1'b1, 1'b0};
4358: data_out = {8'd133, 8'd108, 1'b1, 1'b0};
4359: data_out = {8'd134, 8'd108, 1'b1, 1'b0};
4360: data_out = {8'd135, 8'd108, 1'b1, 1'b0};
4361: data_out = {8'd137, 8'd108, 1'b1, 1'b0};
4362: data_out = {8'd138, 8'd108, 1'b1, 1'b0};
4363: data_out = {8'd139, 8'd108, 1'b1, 1'b0};
4364: data_out = {8'd140, 8'd108, 1'b1, 1'b0};
4365: data_out = {8'd141, 8'd108, 1'b1, 1'b0};
4366: data_out = {8'd143, 8'd108, 1'b1, 1'b0};
4367: data_out = {8'd146, 8'd108, 1'b1, 1'b0};
4368: data_out = {8'd149, 8'd108, 1'b1, 1'b0};
4369: data_out = {8'd54, 8'd113, 1'b1, 1'b0};
4370: data_out = {8'd48, 8'd114, 1'b1, 1'b0};
4371: data_out = {8'd54, 8'd114, 1'b1, 1'b0};
4372: data_out = {8'd81, 8'd114, 1'b1, 1'b0};
4373: data_out = {8'd6, 8'd115, 1'b1, 1'b0};
4374: data_out = {8'd7, 8'd115, 1'b1, 1'b0};
4375: data_out = {8'd8, 8'd115, 1'b1, 1'b0};
4376: data_out = {8'd9, 8'd115, 1'b1, 1'b0};
4377: data_out = {8'd10, 8'd115, 1'b1, 1'b0};
4378: data_out = {8'd13, 8'd115, 1'b1, 1'b0};
4379: data_out = {8'd14, 8'd115, 1'b1, 1'b0};
4380: data_out = {8'd15, 8'd115, 1'b1, 1'b0};
4381: data_out = {8'd16, 8'd115, 1'b1, 1'b0};
4382: data_out = {8'd17, 8'd115, 1'b1, 1'b0};
4383: data_out = {8'd20, 8'd115, 1'b1, 1'b0};
4384: data_out = {8'd21, 8'd115, 1'b1, 1'b0};
4385: data_out = {8'd22, 8'd115, 1'b1, 1'b0};
4386: data_out = {8'd23, 8'd115, 1'b1, 1'b0};
4387: data_out = {8'd24, 8'd115, 1'b1, 1'b0};
4388: data_out = {8'd26, 8'd115, 1'b1, 1'b0};
4389: data_out = {8'd27, 8'd115, 1'b1, 1'b0};
4390: data_out = {8'd28, 8'd115, 1'b1, 1'b0};
4391: data_out = {8'd29, 8'd115, 1'b1, 1'b0};
4392: data_out = {8'd30, 8'd115, 1'b1, 1'b0};
4393: data_out = {8'd31, 8'd115, 1'b1, 1'b0};
4394: data_out = {8'd32, 8'd115, 1'b1, 1'b0};
4395: data_out = {8'd35, 8'd115, 1'b1, 1'b0};
4396: data_out = {8'd39, 8'd115, 1'b1, 1'b0};
4397: data_out = {8'd47, 8'd115, 1'b1, 1'b0};
4398: data_out = {8'd48, 8'd115, 1'b1, 1'b0};
4399: data_out = {8'd49, 8'd115, 1'b1, 1'b0};
4400: data_out = {8'd50, 8'd115, 1'b1, 1'b0};
4401: data_out = {8'd51, 8'd115, 1'b1, 1'b0};
4402: data_out = {8'd54, 8'd115, 1'b1, 1'b0};
4403: data_out = {8'd55, 8'd115, 1'b1, 1'b0};
4404: data_out = {8'd56, 8'd115, 1'b1, 1'b0};
4405: data_out = {8'd57, 8'd115, 1'b1, 1'b0};
4406: data_out = {8'd58, 8'd115, 1'b1, 1'b0};
4407: data_out = {8'd62, 8'd115, 1'b1, 1'b0};
4408: data_out = {8'd63, 8'd115, 1'b1, 1'b0};
4409: data_out = {8'd64, 8'd115, 1'b1, 1'b0};
4410: data_out = {8'd67, 8'd115, 1'b1, 1'b0};
4411: data_out = {8'd68, 8'd115, 1'b1, 1'b0};
4412: data_out = {8'd69, 8'd115, 1'b1, 1'b0};
4413: data_out = {8'd70, 8'd115, 1'b1, 1'b0};
4414: data_out = {8'd71, 8'd115, 1'b1, 1'b0};
4415: data_out = {8'd74, 8'd115, 1'b1, 1'b0};
4416: data_out = {8'd75, 8'd115, 1'b1, 1'b0};
4417: data_out = {8'd76, 8'd115, 1'b1, 1'b0};
4418: data_out = {8'd77, 8'd115, 1'b1, 1'b0};
4419: data_out = {8'd78, 8'd115, 1'b1, 1'b0};
4420: data_out = {8'd80, 8'd115, 1'b1, 1'b0};
4421: data_out = {8'd81, 8'd115, 1'b1, 1'b0};
4422: data_out = {8'd82, 8'd115, 1'b1, 1'b0};
4423: data_out = {8'd83, 8'd115, 1'b1, 1'b0};
4424: data_out = {8'd84, 8'd115, 1'b1, 1'b0};
4425: data_out = {8'd87, 8'd115, 1'b1, 1'b0};
4426: data_out = {8'd88, 8'd115, 1'b1, 1'b0};
4427: data_out = {8'd89, 8'd115, 1'b1, 1'b0};
4428: data_out = {8'd90, 8'd115, 1'b1, 1'b0};
4429: data_out = {8'd91, 8'd115, 1'b1, 1'b0};
4430: data_out = {8'd6, 8'd116, 1'b1, 1'b0};
4431: data_out = {8'd10, 8'd116, 1'b1, 1'b0};
4432: data_out = {8'd13, 8'd116, 1'b1, 1'b0};
4433: data_out = {8'd17, 8'd116, 1'b1, 1'b0};
4434: data_out = {8'd20, 8'd116, 1'b1, 1'b0};
4435: data_out = {8'd24, 8'd116, 1'b1, 1'b0};
4436: data_out = {8'd26, 8'd116, 1'b1, 1'b0};
4437: data_out = {8'd29, 8'd116, 1'b1, 1'b0};
4438: data_out = {8'd32, 8'd116, 1'b1, 1'b0};
4439: data_out = {8'd35, 8'd116, 1'b1, 1'b0};
4440: data_out = {8'd39, 8'd116, 1'b1, 1'b0};
4441: data_out = {8'd48, 8'd116, 1'b1, 1'b0};
4442: data_out = {8'd54, 8'd116, 1'b1, 1'b0};
4443: data_out = {8'd58, 8'd116, 1'b1, 1'b0};
4444: data_out = {8'd62, 8'd116, 1'b1, 1'b0};
4445: data_out = {8'd64, 8'd116, 1'b1, 1'b0};
4446: data_out = {8'd67, 8'd116, 1'b1, 1'b0};
4447: data_out = {8'd71, 8'd116, 1'b1, 1'b0};
4448: data_out = {8'd74, 8'd116, 1'b1, 1'b0};
4449: data_out = {8'd78, 8'd116, 1'b1, 1'b0};
4450: data_out = {8'd81, 8'd116, 1'b1, 1'b0};
4451: data_out = {8'd87, 8'd116, 1'b1, 1'b0};
4452: data_out = {8'd91, 8'd116, 1'b1, 1'b0};
4453: data_out = {8'd6, 8'd117, 1'b1, 1'b0};
4454: data_out = {8'd10, 8'd117, 1'b1, 1'b0};
4455: data_out = {8'd13, 8'd117, 1'b1, 1'b0};
4456: data_out = {8'd17, 8'd117, 1'b1, 1'b0};
4457: data_out = {8'd20, 8'd117, 1'b1, 1'b0};
4458: data_out = {8'd24, 8'd117, 1'b1, 1'b0};
4459: data_out = {8'd26, 8'd117, 1'b1, 1'b0};
4460: data_out = {8'd29, 8'd117, 1'b1, 1'b0};
4461: data_out = {8'd32, 8'd117, 1'b1, 1'b0};
4462: data_out = {8'd35, 8'd117, 1'b1, 1'b0};
4463: data_out = {8'd39, 8'd117, 1'b1, 1'b0};
4464: data_out = {8'd48, 8'd117, 1'b1, 1'b0};
4465: data_out = {8'd54, 8'd117, 1'b1, 1'b0};
4466: data_out = {8'd58, 8'd117, 1'b1, 1'b0};
4467: data_out = {8'd62, 8'd117, 1'b1, 1'b0};
4468: data_out = {8'd67, 8'd117, 1'b1, 1'b0};
4469: data_out = {8'd71, 8'd117, 1'b1, 1'b0};
4470: data_out = {8'd78, 8'd117, 1'b1, 1'b0};
4471: data_out = {8'd81, 8'd117, 1'b1, 1'b0};
4472: data_out = {8'd87, 8'd117, 1'b1, 1'b0};
4473: data_out = {8'd6, 8'd118, 1'b1, 1'b0};
4474: data_out = {8'd7, 8'd118, 1'b1, 1'b0};
4475: data_out = {8'd8, 8'd118, 1'b1, 1'b0};
4476: data_out = {8'd9, 8'd118, 1'b1, 1'b0};
4477: data_out = {8'd13, 8'd118, 1'b1, 1'b0};
4478: data_out = {8'd17, 8'd118, 1'b1, 1'b0};
4479: data_out = {8'd20, 8'd118, 1'b1, 1'b0};
4480: data_out = {8'd21, 8'd118, 1'b1, 1'b0};
4481: data_out = {8'd22, 8'd118, 1'b1, 1'b0};
4482: data_out = {8'd23, 8'd118, 1'b1, 1'b0};
4483: data_out = {8'd26, 8'd118, 1'b1, 1'b0};
4484: data_out = {8'd29, 8'd118, 1'b1, 1'b0};
4485: data_out = {8'd32, 8'd118, 1'b1, 1'b0};
4486: data_out = {8'd35, 8'd118, 1'b1, 1'b0};
4487: data_out = {8'd39, 8'd118, 1'b1, 1'b0};
4488: data_out = {8'd48, 8'd118, 1'b1, 1'b0};
4489: data_out = {8'd54, 8'd118, 1'b1, 1'b0};
4490: data_out = {8'd58, 8'd118, 1'b1, 1'b0};
4491: data_out = {8'd62, 8'd118, 1'b1, 1'b0};
4492: data_out = {8'd67, 8'd118, 1'b1, 1'b0};
4493: data_out = {8'd68, 8'd118, 1'b1, 1'b0};
4494: data_out = {8'd69, 8'd118, 1'b1, 1'b0};
4495: data_out = {8'd70, 8'd118, 1'b1, 1'b0};
4496: data_out = {8'd75, 8'd118, 1'b1, 1'b0};
4497: data_out = {8'd76, 8'd118, 1'b1, 1'b0};
4498: data_out = {8'd77, 8'd118, 1'b1, 1'b0};
4499: data_out = {8'd78, 8'd118, 1'b1, 1'b0};
4500: data_out = {8'd81, 8'd118, 1'b1, 1'b0};
4501: data_out = {8'd87, 8'd118, 1'b1, 1'b0};
4502: data_out = {8'd88, 8'd118, 1'b1, 1'b0};
4503: data_out = {8'd89, 8'd118, 1'b1, 1'b0};
4504: data_out = {8'd90, 8'd118, 1'b1, 1'b0};
4505: data_out = {8'd91, 8'd118, 1'b1, 1'b0};
4506: data_out = {8'd6, 8'd119, 1'b1, 1'b0};
4507: data_out = {8'd13, 8'd119, 1'b1, 1'b0};
4508: data_out = {8'd17, 8'd119, 1'b1, 1'b0};
4509: data_out = {8'd20, 8'd119, 1'b1, 1'b0};
4510: data_out = {8'd26, 8'd119, 1'b1, 1'b0};
4511: data_out = {8'd29, 8'd119, 1'b1, 1'b0};
4512: data_out = {8'd32, 8'd119, 1'b1, 1'b0};
4513: data_out = {8'd35, 8'd119, 1'b1, 1'b0};
4514: data_out = {8'd39, 8'd119, 1'b1, 1'b0};
4515: data_out = {8'd48, 8'd119, 1'b1, 1'b0};
4516: data_out = {8'd54, 8'd119, 1'b1, 1'b0};
4517: data_out = {8'd58, 8'd119, 1'b1, 1'b0};
4518: data_out = {8'd62, 8'd119, 1'b1, 1'b0};
4519: data_out = {8'd67, 8'd119, 1'b1, 1'b0};
4520: data_out = {8'd74, 8'd119, 1'b1, 1'b0};
4521: data_out = {8'd78, 8'd119, 1'b1, 1'b0};
4522: data_out = {8'd81, 8'd119, 1'b1, 1'b0};
4523: data_out = {8'd91, 8'd119, 1'b1, 1'b0};
4524: data_out = {8'd6, 8'd120, 1'b1, 1'b0};
4525: data_out = {8'd13, 8'd120, 1'b1, 1'b0};
4526: data_out = {8'd17, 8'd120, 1'b1, 1'b0};
4527: data_out = {8'd20, 8'd120, 1'b1, 1'b0};
4528: data_out = {8'd26, 8'd120, 1'b1, 1'b0};
4529: data_out = {8'd29, 8'd120, 1'b1, 1'b0};
4530: data_out = {8'd32, 8'd120, 1'b1, 1'b0};
4531: data_out = {8'd35, 8'd120, 1'b1, 1'b0};
4532: data_out = {8'd39, 8'd120, 1'b1, 1'b0};
4533: data_out = {8'd48, 8'd120, 1'b1, 1'b0};
4534: data_out = {8'd54, 8'd120, 1'b1, 1'b0};
4535: data_out = {8'd58, 8'd120, 1'b1, 1'b0};
4536: data_out = {8'd62, 8'd120, 1'b1, 1'b0};
4537: data_out = {8'd67, 8'd120, 1'b1, 1'b0};
4538: data_out = {8'd74, 8'd120, 1'b1, 1'b0};
4539: data_out = {8'd78, 8'd120, 1'b1, 1'b0};
4540: data_out = {8'd81, 8'd120, 1'b1, 1'b0};
4541: data_out = {8'd91, 8'd120, 1'b1, 1'b0};
4542: data_out = {8'd6, 8'd121, 1'b1, 1'b0};
4543: data_out = {8'd7, 8'd121, 1'b1, 1'b0};
4544: data_out = {8'd8, 8'd121, 1'b1, 1'b0};
4545: data_out = {8'd9, 8'd121, 1'b1, 1'b0};
4546: data_out = {8'd10, 8'd121, 1'b1, 1'b0};
4547: data_out = {8'd13, 8'd121, 1'b1, 1'b0};
4548: data_out = {8'd17, 8'd121, 1'b1, 1'b0};
4549: data_out = {8'd20, 8'd121, 1'b1, 1'b0};
4550: data_out = {8'd21, 8'd121, 1'b1, 1'b0};
4551: data_out = {8'd22, 8'd121, 1'b1, 1'b0};
4552: data_out = {8'd23, 8'd121, 1'b1, 1'b0};
4553: data_out = {8'd24, 8'd121, 1'b1, 1'b0};
4554: data_out = {8'd26, 8'd121, 1'b1, 1'b0};
4555: data_out = {8'd29, 8'd121, 1'b1, 1'b0};
4556: data_out = {8'd32, 8'd121, 1'b1, 1'b0};
4557: data_out = {8'd35, 8'd121, 1'b1, 1'b0};
4558: data_out = {8'd36, 8'd121, 1'b1, 1'b0};
4559: data_out = {8'd37, 8'd121, 1'b1, 1'b0};
4560: data_out = {8'd38, 8'd121, 1'b1, 1'b0};
4561: data_out = {8'd39, 8'd121, 1'b1, 1'b0};
4562: data_out = {8'd48, 8'd121, 1'b1, 1'b0};
4563: data_out = {8'd49, 8'd121, 1'b1, 1'b0};
4564: data_out = {8'd50, 8'd121, 1'b1, 1'b0};
4565: data_out = {8'd51, 8'd121, 1'b1, 1'b0};
4566: data_out = {8'd52, 8'd121, 1'b1, 1'b0};
4567: data_out = {8'd54, 8'd121, 1'b1, 1'b0};
4568: data_out = {8'd58, 8'd121, 1'b1, 1'b0};
4569: data_out = {8'd60, 8'd121, 1'b1, 1'b0};
4570: data_out = {8'd61, 8'd121, 1'b1, 1'b0};
4571: data_out = {8'd62, 8'd121, 1'b1, 1'b0};
4572: data_out = {8'd63, 8'd121, 1'b1, 1'b0};
4573: data_out = {8'd64, 8'd121, 1'b1, 1'b0};
4574: data_out = {8'd65, 8'd121, 1'b1, 1'b0};
4575: data_out = {8'd67, 8'd121, 1'b1, 1'b0};
4576: data_out = {8'd68, 8'd121, 1'b1, 1'b0};
4577: data_out = {8'd69, 8'd121, 1'b1, 1'b0};
4578: data_out = {8'd70, 8'd121, 1'b1, 1'b0};
4579: data_out = {8'd71, 8'd121, 1'b1, 1'b0};
4580: data_out = {8'd74, 8'd121, 1'b1, 1'b0};
4581: data_out = {8'd75, 8'd121, 1'b1, 1'b0};
4582: data_out = {8'd76, 8'd121, 1'b1, 1'b0};
4583: data_out = {8'd77, 8'd121, 1'b1, 1'b0};
4584: data_out = {8'd78, 8'd121, 1'b1, 1'b0};
4585: data_out = {8'd81, 8'd121, 1'b1, 1'b0};
4586: data_out = {8'd82, 8'd121, 1'b1, 1'b0};
4587: data_out = {8'd83, 8'd121, 1'b1, 1'b0};
4588: data_out = {8'd84, 8'd121, 1'b1, 1'b0};
4589: data_out = {8'd85, 8'd121, 1'b1, 1'b0};
4590: data_out = {8'd87, 8'd121, 1'b1, 1'b0};
4591: data_out = {8'd88, 8'd121, 1'b1, 1'b0};
4592: data_out = {8'd89, 8'd121, 1'b1, 1'b0};
4593: data_out = {8'd90, 8'd121, 1'b1, 1'b0};
4594: data_out = {8'd91, 8'd121, 1'b1, 1'b0};
4595: data_out = {8'd95, 8'd121, 1'b1, 1'b0};
4596: data_out = {8'd39, 8'd122, 1'b1, 1'b0};
4597: data_out = {8'd39, 8'd123, 1'b1, 1'b0};
4598: data_out = {8'd35, 8'd124, 1'b1, 1'b0};
4599: data_out = {8'd36, 8'd124, 1'b1, 1'b0};
4600: data_out = {8'd37, 8'd124, 1'b1, 1'b0};
4601: data_out = {8'd38, 8'd124, 1'b1, 1'b0};
4602: data_out = {8'd39, 8'd124, 1'b1, 1'b0};
4603: data_out = {8'd7, 8'd138, 1'b1, 1'b0};
4604: data_out = {8'd8, 8'd138, 1'b1, 1'b0};
4605: data_out = {8'd9, 8'd138, 1'b1, 1'b0};
4606: data_out = {8'd10, 8'd138, 1'b1, 1'b0};
4607: data_out = {8'd7, 8'd139, 1'b1, 1'b0};
4608: data_out = {8'd10, 8'd139, 1'b1, 1'b0};
4609: data_out = {8'd13, 8'd139, 1'b1, 1'b0};
4610: data_out = {8'd14, 8'd139, 1'b1, 1'b0};
4611: data_out = {8'd15, 8'd139, 1'b1, 1'b0};
4612: data_out = {8'd21, 8'd139, 1'b1, 1'b0};
4613: data_out = {8'd7, 8'd140, 1'b1, 1'b0};
4614: data_out = {8'd15, 8'd140, 1'b1, 1'b0};
4615: data_out = {8'd5, 8'd141, 1'b1, 1'b0};
4616: data_out = {8'd6, 8'd141, 1'b1, 1'b0};
4617: data_out = {8'd7, 8'd141, 1'b1, 1'b0};
4618: data_out = {8'd8, 8'd141, 1'b1, 1'b0};
4619: data_out = {8'd9, 8'd141, 1'b1, 1'b0};
4620: data_out = {8'd10, 8'd141, 1'b1, 1'b0};
4621: data_out = {8'd15, 8'd141, 1'b1, 1'b0};
4622: data_out = {8'd19, 8'd141, 1'b1, 1'b0};
4623: data_out = {8'd20, 8'd141, 1'b1, 1'b0};
4624: data_out = {8'd21, 8'd141, 1'b1, 1'b0};
4625: data_out = {8'd25, 8'd141, 1'b1, 1'b0};
4626: data_out = {8'd26, 8'd141, 1'b1, 1'b0};
4627: data_out = {8'd27, 8'd141, 1'b1, 1'b0};
4628: data_out = {8'd28, 8'd141, 1'b1, 1'b0};
4629: data_out = {8'd29, 8'd141, 1'b1, 1'b0};
4630: data_out = {8'd38, 8'd141, 1'b1, 1'b0};
4631: data_out = {8'd39, 8'd141, 1'b1, 1'b0};
4632: data_out = {8'd40, 8'd141, 1'b1, 1'b0};
4633: data_out = {8'd41, 8'd141, 1'b1, 1'b0};
4634: data_out = {8'd42, 8'd141, 1'b1, 1'b0};
4635: data_out = {8'd44, 8'd141, 1'b1, 1'b0};
4636: data_out = {8'd49, 8'd141, 1'b1, 1'b0};
4637: data_out = {8'd53, 8'd141, 1'b1, 1'b0};
4638: data_out = {8'd54, 8'd141, 1'b1, 1'b0};
4639: data_out = {8'd58, 8'd141, 1'b1, 1'b0};
4640: data_out = {8'd59, 8'd141, 1'b1, 1'b0};
4641: data_out = {8'd60, 8'd141, 1'b1, 1'b0};
4642: data_out = {8'd61, 8'd141, 1'b1, 1'b0};
4643: data_out = {8'd62, 8'd141, 1'b1, 1'b0};
4644: data_out = {8'd77, 8'd141, 1'b1, 1'b0};
4645: data_out = {8'd78, 8'd141, 1'b1, 1'b0};
4646: data_out = {8'd79, 8'd141, 1'b1, 1'b0};
4647: data_out = {8'd80, 8'd141, 1'b1, 1'b0};
4648: data_out = {8'd81, 8'd141, 1'b1, 1'b0};
4649: data_out = {8'd83, 8'd141, 1'b1, 1'b0};
4650: data_out = {8'd88, 8'd141, 1'b1, 1'b0};
4651: data_out = {8'd92, 8'd141, 1'b1, 1'b0};
4652: data_out = {8'd93, 8'd141, 1'b1, 1'b0};
4653: data_out = {8'd98, 8'd141, 1'b1, 1'b0};
4654: data_out = {8'd99, 8'd141, 1'b1, 1'b0};
4655: data_out = {8'd100, 8'd141, 1'b1, 1'b0};
4656: data_out = {8'd115, 8'd141, 1'b1, 1'b0};
4657: data_out = {8'd116, 8'd141, 1'b1, 1'b0};
4658: data_out = {8'd117, 8'd141, 1'b1, 1'b0};
4659: data_out = {8'd118, 8'd141, 1'b1, 1'b0};
4660: data_out = {8'd119, 8'd141, 1'b1, 1'b0};
4661: data_out = {8'd121, 8'd141, 1'b1, 1'b0};
4662: data_out = {8'd126, 8'd141, 1'b1, 1'b0};
4663: data_out = {8'd130, 8'd141, 1'b1, 1'b0};
4664: data_out = {8'd131, 8'd141, 1'b1, 1'b0};
4665: data_out = {8'd135, 8'd141, 1'b1, 1'b0};
4666: data_out = {8'd136, 8'd141, 1'b1, 1'b0};
4667: data_out = {8'd137, 8'd141, 1'b1, 1'b0};
4668: data_out = {8'd138, 8'd141, 1'b1, 1'b0};
4669: data_out = {8'd153, 8'd141, 1'b1, 1'b0};
4670: data_out = {8'd154, 8'd141, 1'b1, 1'b0};
4671: data_out = {8'd155, 8'd141, 1'b1, 1'b0};
4672: data_out = {8'd156, 8'd141, 1'b1, 1'b0};
4673: data_out = {8'd157, 8'd141, 1'b1, 1'b0};
4674: data_out = {8'd159, 8'd141, 1'b1, 1'b0};
4675: data_out = {8'd164, 8'd141, 1'b1, 1'b0};
4676: data_out = {8'd168, 8'd141, 1'b1, 1'b0};
4677: data_out = {8'd169, 8'd141, 1'b1, 1'b0};
4678: data_out = {8'd173, 8'd141, 1'b1, 1'b0};
4679: data_out = {8'd174, 8'd141, 1'b1, 1'b0};
4680: data_out = {8'd175, 8'd141, 1'b1, 1'b0};
4681: data_out = {8'd176, 8'd141, 1'b1, 1'b0};
4682: data_out = {8'd177, 8'd141, 1'b1, 1'b0};
4683: data_out = {8'd186, 8'd141, 1'b1, 1'b0};
4684: data_out = {8'd190, 8'd141, 1'b1, 1'b0};
4685: data_out = {8'd193, 8'd141, 1'b1, 1'b0};
4686: data_out = {8'd194, 8'd141, 1'b1, 1'b0};
4687: data_out = {8'd195, 8'd141, 1'b1, 1'b0};
4688: data_out = {8'd196, 8'd141, 1'b1, 1'b0};
4689: data_out = {8'd197, 8'd141, 1'b1, 1'b0};
4690: data_out = {8'd7, 8'd142, 1'b1, 1'b0};
4691: data_out = {8'd15, 8'd142, 1'b1, 1'b0};
4692: data_out = {8'd21, 8'd142, 1'b1, 1'b0};
4693: data_out = {8'd25, 8'd142, 1'b1, 1'b0};
4694: data_out = {8'd29, 8'd142, 1'b1, 1'b0};
4695: data_out = {8'd38, 8'd142, 1'b1, 1'b0};
4696: data_out = {8'd42, 8'd142, 1'b1, 1'b0};
4697: data_out = {8'd44, 8'd142, 1'b1, 1'b0};
4698: data_out = {8'd49, 8'd142, 1'b1, 1'b0};
4699: data_out = {8'd52, 8'd142, 1'b1, 1'b0};
4700: data_out = {8'd54, 8'd142, 1'b1, 1'b0};
4701: data_out = {8'd58, 8'd142, 1'b1, 1'b0};
4702: data_out = {8'd77, 8'd142, 1'b1, 1'b0};
4703: data_out = {8'd81, 8'd142, 1'b1, 1'b0};
4704: data_out = {8'd83, 8'd142, 1'b1, 1'b0};
4705: data_out = {8'd88, 8'd142, 1'b1, 1'b0};
4706: data_out = {8'd91, 8'd142, 1'b1, 1'b0};
4707: data_out = {8'd93, 8'd142, 1'b1, 1'b0};
4708: data_out = {8'd98, 8'd142, 1'b1, 1'b0};
4709: data_out = {8'd100, 8'd142, 1'b1, 1'b0};
4710: data_out = {8'd115, 8'd142, 1'b1, 1'b0};
4711: data_out = {8'd119, 8'd142, 1'b1, 1'b0};
4712: data_out = {8'd121, 8'd142, 1'b1, 1'b0};
4713: data_out = {8'd126, 8'd142, 1'b1, 1'b0};
4714: data_out = {8'd129, 8'd142, 1'b1, 1'b0};
4715: data_out = {8'd131, 8'd142, 1'b1, 1'b0};
4716: data_out = {8'd135, 8'd142, 1'b1, 1'b0};
4717: data_out = {8'd138, 8'd142, 1'b1, 1'b0};
4718: data_out = {8'd153, 8'd142, 1'b1, 1'b0};
4719: data_out = {8'd157, 8'd142, 1'b1, 1'b0};
4720: data_out = {8'd159, 8'd142, 1'b1, 1'b0};
4721: data_out = {8'd164, 8'd142, 1'b1, 1'b0};
4722: data_out = {8'd167, 8'd142, 1'b1, 1'b0};
4723: data_out = {8'd169, 8'd142, 1'b1, 1'b0};
4724: data_out = {8'd173, 8'd142, 1'b1, 1'b0};
4725: data_out = {8'd177, 8'd142, 1'b1, 1'b0};
4726: data_out = {8'd186, 8'd142, 1'b1, 1'b0};
4727: data_out = {8'd190, 8'd142, 1'b1, 1'b0};
4728: data_out = {8'd193, 8'd142, 1'b1, 1'b0};
4729: data_out = {8'd197, 8'd142, 1'b1, 1'b0};
4730: data_out = {8'd7, 8'd143, 1'b1, 1'b0};
4731: data_out = {8'd15, 8'd143, 1'b1, 1'b0};
4732: data_out = {8'd21, 8'd143, 1'b1, 1'b0};
4733: data_out = {8'd25, 8'd143, 1'b1, 1'b0};
4734: data_out = {8'd29, 8'd143, 1'b1, 1'b0};
4735: data_out = {8'd38, 8'd143, 1'b1, 1'b0};
4736: data_out = {8'd44, 8'd143, 1'b1, 1'b0};
4737: data_out = {8'd49, 8'd143, 1'b1, 1'b0};
4738: data_out = {8'd54, 8'd143, 1'b1, 1'b0};
4739: data_out = {8'd58, 8'd143, 1'b1, 1'b0};
4740: data_out = {8'd77, 8'd143, 1'b1, 1'b0};
4741: data_out = {8'd83, 8'd143, 1'b1, 1'b0};
4742: data_out = {8'd88, 8'd143, 1'b1, 1'b0};
4743: data_out = {8'd93, 8'd143, 1'b1, 1'b0};
4744: data_out = {8'd97, 8'd143, 1'b1, 1'b0};
4745: data_out = {8'd100, 8'd143, 1'b1, 1'b0};
4746: data_out = {8'd115, 8'd143, 1'b1, 1'b0};
4747: data_out = {8'd121, 8'd143, 1'b1, 1'b0};
4748: data_out = {8'd126, 8'd143, 1'b1, 1'b0};
4749: data_out = {8'd131, 8'd143, 1'b1, 1'b0};
4750: data_out = {8'd137, 8'd143, 1'b1, 1'b0};
4751: data_out = {8'd153, 8'd143, 1'b1, 1'b0};
4752: data_out = {8'd159, 8'd143, 1'b1, 1'b0};
4753: data_out = {8'd164, 8'd143, 1'b1, 1'b0};
4754: data_out = {8'd169, 8'd143, 1'b1, 1'b0};
4755: data_out = {8'd177, 8'd143, 1'b1, 1'b0};
4756: data_out = {8'd186, 8'd143, 1'b1, 1'b0};
4757: data_out = {8'd190, 8'd143, 1'b1, 1'b0};
4758: data_out = {8'd193, 8'd143, 1'b1, 1'b0};
4759: data_out = {8'd197, 8'd143, 1'b1, 1'b0};
4760: data_out = {8'd7, 8'd144, 1'b1, 1'b0};
4761: data_out = {8'd15, 8'd144, 1'b1, 1'b0};
4762: data_out = {8'd21, 8'd144, 1'b1, 1'b0};
4763: data_out = {8'd25, 8'd144, 1'b1, 1'b0};
4764: data_out = {8'd29, 8'd144, 1'b1, 1'b0};
4765: data_out = {8'd38, 8'd144, 1'b1, 1'b0};
4766: data_out = {8'd39, 8'd144, 1'b1, 1'b0};
4767: data_out = {8'd40, 8'd144, 1'b1, 1'b0};
4768: data_out = {8'd41, 8'd144, 1'b1, 1'b0};
4769: data_out = {8'd42, 8'd144, 1'b1, 1'b0};
4770: data_out = {8'd44, 8'd144, 1'b1, 1'b0};
4771: data_out = {8'd46, 8'd144, 1'b1, 1'b0};
4772: data_out = {8'd49, 8'd144, 1'b1, 1'b0};
4773: data_out = {8'd54, 8'd144, 1'b1, 1'b0};
4774: data_out = {8'd58, 8'd144, 1'b1, 1'b0};
4775: data_out = {8'd59, 8'd144, 1'b1, 1'b0};
4776: data_out = {8'd60, 8'd144, 1'b1, 1'b0};
4777: data_out = {8'd61, 8'd144, 1'b1, 1'b0};
4778: data_out = {8'd62, 8'd144, 1'b1, 1'b0};
4779: data_out = {8'd77, 8'd144, 1'b1, 1'b0};
4780: data_out = {8'd78, 8'd144, 1'b1, 1'b0};
4781: data_out = {8'd79, 8'd144, 1'b1, 1'b0};
4782: data_out = {8'd80, 8'd144, 1'b1, 1'b0};
4783: data_out = {8'd81, 8'd144, 1'b1, 1'b0};
4784: data_out = {8'd83, 8'd144, 1'b1, 1'b0};
4785: data_out = {8'd85, 8'd144, 1'b1, 1'b0};
4786: data_out = {8'd88, 8'd144, 1'b1, 1'b0};
4787: data_out = {8'd93, 8'd144, 1'b1, 1'b0};
4788: data_out = {8'd96, 8'd144, 1'b1, 1'b0};
4789: data_out = {8'd100, 8'd144, 1'b1, 1'b0};
4790: data_out = {8'd115, 8'd144, 1'b1, 1'b0};
4791: data_out = {8'd116, 8'd144, 1'b1, 1'b0};
4792: data_out = {8'd117, 8'd144, 1'b1, 1'b0};
4793: data_out = {8'd118, 8'd144, 1'b1, 1'b0};
4794: data_out = {8'd119, 8'd144, 1'b1, 1'b0};
4795: data_out = {8'd121, 8'd144, 1'b1, 1'b0};
4796: data_out = {8'd123, 8'd144, 1'b1, 1'b0};
4797: data_out = {8'd126, 8'd144, 1'b1, 1'b0};
4798: data_out = {8'd131, 8'd144, 1'b1, 1'b0};
4799: data_out = {8'd136, 8'd144, 1'b1, 1'b0};
4800: data_out = {8'd137, 8'd144, 1'b1, 1'b0};
4801: data_out = {8'd138, 8'd144, 1'b1, 1'b0};
4802: data_out = {8'd153, 8'd144, 1'b1, 1'b0};
4803: data_out = {8'd154, 8'd144, 1'b1, 1'b0};
4804: data_out = {8'd155, 8'd144, 1'b1, 1'b0};
4805: data_out = {8'd156, 8'd144, 1'b1, 1'b0};
4806: data_out = {8'd157, 8'd144, 1'b1, 1'b0};
4807: data_out = {8'd159, 8'd144, 1'b1, 1'b0};
4808: data_out = {8'd161, 8'd144, 1'b1, 1'b0};
4809: data_out = {8'd164, 8'd144, 1'b1, 1'b0};
4810: data_out = {8'd169, 8'd144, 1'b1, 1'b0};
4811: data_out = {8'd173, 8'd144, 1'b1, 1'b0};
4812: data_out = {8'd174, 8'd144, 1'b1, 1'b0};
4813: data_out = {8'd175, 8'd144, 1'b1, 1'b0};
4814: data_out = {8'd176, 8'd144, 1'b1, 1'b0};
4815: data_out = {8'd177, 8'd144, 1'b1, 1'b0};
4816: data_out = {8'd186, 8'd144, 1'b1, 1'b0};
4817: data_out = {8'd190, 8'd144, 1'b1, 1'b0};
4818: data_out = {8'd193, 8'd144, 1'b1, 1'b0};
4819: data_out = {8'd197, 8'd144, 1'b1, 1'b0};
4820: data_out = {8'd7, 8'd145, 1'b1, 1'b0};
4821: data_out = {8'd15, 8'd145, 1'b1, 1'b0};
4822: data_out = {8'd21, 8'd145, 1'b1, 1'b0};
4823: data_out = {8'd25, 8'd145, 1'b1, 1'b0};
4824: data_out = {8'd29, 8'd145, 1'b1, 1'b0};
4825: data_out = {8'd42, 8'd145, 1'b1, 1'b0};
4826: data_out = {8'd44, 8'd145, 1'b1, 1'b0};
4827: data_out = {8'd46, 8'd145, 1'b1, 1'b0};
4828: data_out = {8'd47, 8'd145, 1'b1, 1'b0};
4829: data_out = {8'd49, 8'd145, 1'b1, 1'b0};
4830: data_out = {8'd54, 8'd145, 1'b1, 1'b0};
4831: data_out = {8'd58, 8'd145, 1'b1, 1'b0};
4832: data_out = {8'd62, 8'd145, 1'b1, 1'b0};
4833: data_out = {8'd81, 8'd145, 1'b1, 1'b0};
4834: data_out = {8'd83, 8'd145, 1'b1, 1'b0};
4835: data_out = {8'd85, 8'd145, 1'b1, 1'b0};
4836: data_out = {8'd86, 8'd145, 1'b1, 1'b0};
4837: data_out = {8'd88, 8'd145, 1'b1, 1'b0};
4838: data_out = {8'd93, 8'd145, 1'b1, 1'b0};
4839: data_out = {8'd96, 8'd145, 1'b1, 1'b0};
4840: data_out = {8'd97, 8'd145, 1'b1, 1'b0};
4841: data_out = {8'd98, 8'd145, 1'b1, 1'b0};
4842: data_out = {8'd99, 8'd145, 1'b1, 1'b0};
4843: data_out = {8'd100, 8'd145, 1'b1, 1'b0};
4844: data_out = {8'd101, 8'd145, 1'b1, 1'b0};
4845: data_out = {8'd119, 8'd145, 1'b1, 1'b0};
4846: data_out = {8'd121, 8'd145, 1'b1, 1'b0};
4847: data_out = {8'd123, 8'd145, 1'b1, 1'b0};
4848: data_out = {8'd124, 8'd145, 1'b1, 1'b0};
4849: data_out = {8'd126, 8'd145, 1'b1, 1'b0};
4850: data_out = {8'd131, 8'd145, 1'b1, 1'b0};
4851: data_out = {8'd138, 8'd145, 1'b1, 1'b0};
4852: data_out = {8'd157, 8'd145, 1'b1, 1'b0};
4853: data_out = {8'd159, 8'd145, 1'b1, 1'b0};
4854: data_out = {8'd161, 8'd145, 1'b1, 1'b0};
4855: data_out = {8'd162, 8'd145, 1'b1, 1'b0};
4856: data_out = {8'd164, 8'd145, 1'b1, 1'b0};
4857: data_out = {8'd169, 8'd145, 1'b1, 1'b0};
4858: data_out = {8'd173, 8'd145, 1'b1, 1'b0};
4859: data_out = {8'd186, 8'd145, 1'b1, 1'b0};
4860: data_out = {8'd190, 8'd145, 1'b1, 1'b0};
4861: data_out = {8'd193, 8'd145, 1'b1, 1'b0};
4862: data_out = {8'd197, 8'd145, 1'b1, 1'b0};
4863: data_out = {8'd7, 8'd146, 1'b1, 1'b0};
4864: data_out = {8'd15, 8'd146, 1'b1, 1'b0};
4865: data_out = {8'd21, 8'd146, 1'b1, 1'b0};
4866: data_out = {8'd25, 8'd146, 1'b1, 1'b0};
4867: data_out = {8'd29, 8'd146, 1'b1, 1'b0};
4868: data_out = {8'd42, 8'd146, 1'b1, 1'b0};
4869: data_out = {8'd44, 8'd146, 1'b1, 1'b0};
4870: data_out = {8'd45, 8'd146, 1'b1, 1'b0};
4871: data_out = {8'd48, 8'd146, 1'b1, 1'b0};
4872: data_out = {8'd49, 8'd146, 1'b1, 1'b0};
4873: data_out = {8'd54, 8'd146, 1'b1, 1'b0};
4874: data_out = {8'd62, 8'd146, 1'b1, 1'b0};
4875: data_out = {8'd81, 8'd146, 1'b1, 1'b0};
4876: data_out = {8'd83, 8'd146, 1'b1, 1'b0};
4877: data_out = {8'd84, 8'd146, 1'b1, 1'b0};
4878: data_out = {8'd87, 8'd146, 1'b1, 1'b0};
4879: data_out = {8'd88, 8'd146, 1'b1, 1'b0};
4880: data_out = {8'd93, 8'd146, 1'b1, 1'b0};
4881: data_out = {8'd100, 8'd146, 1'b1, 1'b0};
4882: data_out = {8'd119, 8'd146, 1'b1, 1'b0};
4883: data_out = {8'd121, 8'd146, 1'b1, 1'b0};
4884: data_out = {8'd122, 8'd146, 1'b1, 1'b0};
4885: data_out = {8'd125, 8'd146, 1'b1, 1'b0};
4886: data_out = {8'd126, 8'd146, 1'b1, 1'b0};
4887: data_out = {8'd131, 8'd146, 1'b1, 1'b0};
4888: data_out = {8'd138, 8'd146, 1'b1, 1'b0};
4889: data_out = {8'd157, 8'd146, 1'b1, 1'b0};
4890: data_out = {8'd159, 8'd146, 1'b1, 1'b0};
4891: data_out = {8'd160, 8'd146, 1'b1, 1'b0};
4892: data_out = {8'd163, 8'd146, 1'b1, 1'b0};
4893: data_out = {8'd164, 8'd146, 1'b1, 1'b0};
4894: data_out = {8'd169, 8'd146, 1'b1, 1'b0};
4895: data_out = {8'd173, 8'd146, 1'b1, 1'b0};
4896: data_out = {8'd186, 8'd146, 1'b1, 1'b0};
4897: data_out = {8'd190, 8'd146, 1'b1, 1'b0};
4898: data_out = {8'd193, 8'd146, 1'b1, 1'b0};
4899: data_out = {8'd197, 8'd146, 1'b1, 1'b0};
4900: data_out = {8'd5, 8'd147, 1'b1, 1'b0};
4901: data_out = {8'd6, 8'd147, 1'b1, 1'b0};
4902: data_out = {8'd7, 8'd147, 1'b1, 1'b0};
4903: data_out = {8'd8, 8'd147, 1'b1, 1'b0};
4904: data_out = {8'd9, 8'd147, 1'b1, 1'b0};
4905: data_out = {8'd10, 8'd147, 1'b1, 1'b0};
4906: data_out = {8'd13, 8'd147, 1'b1, 1'b0};
4907: data_out = {8'd14, 8'd147, 1'b1, 1'b0};
4908: data_out = {8'd15, 8'd147, 1'b1, 1'b0};
4909: data_out = {8'd16, 8'd147, 1'b1, 1'b0};
4910: data_out = {8'd17, 8'd147, 1'b1, 1'b0};
4911: data_out = {8'd19, 8'd147, 1'b1, 1'b0};
4912: data_out = {8'd20, 8'd147, 1'b1, 1'b0};
4913: data_out = {8'd21, 8'd147, 1'b1, 1'b0};
4914: data_out = {8'd22, 8'd147, 1'b1, 1'b0};
4915: data_out = {8'd23, 8'd147, 1'b1, 1'b0};
4916: data_out = {8'd25, 8'd147, 1'b1, 1'b0};
4917: data_out = {8'd26, 8'd147, 1'b1, 1'b0};
4918: data_out = {8'd27, 8'd147, 1'b1, 1'b0};
4919: data_out = {8'd28, 8'd147, 1'b1, 1'b0};
4920: data_out = {8'd29, 8'd147, 1'b1, 1'b0};
4921: data_out = {8'd38, 8'd147, 1'b1, 1'b0};
4922: data_out = {8'd39, 8'd147, 1'b1, 1'b0};
4923: data_out = {8'd40, 8'd147, 1'b1, 1'b0};
4924: data_out = {8'd41, 8'd147, 1'b1, 1'b0};
4925: data_out = {8'd42, 8'd147, 1'b1, 1'b0};
4926: data_out = {8'd44, 8'd147, 1'b1, 1'b0};
4927: data_out = {8'd49, 8'd147, 1'b1, 1'b0};
4928: data_out = {8'd52, 8'd147, 1'b1, 1'b0};
4929: data_out = {8'd53, 8'd147, 1'b1, 1'b0};
4930: data_out = {8'd54, 8'd147, 1'b1, 1'b0};
4931: data_out = {8'd55, 8'd147, 1'b1, 1'b0};
4932: data_out = {8'd56, 8'd147, 1'b1, 1'b0};
4933: data_out = {8'd58, 8'd147, 1'b1, 1'b0};
4934: data_out = {8'd59, 8'd147, 1'b1, 1'b0};
4935: data_out = {8'd60, 8'd147, 1'b1, 1'b0};
4936: data_out = {8'd61, 8'd147, 1'b1, 1'b0};
4937: data_out = {8'd62, 8'd147, 1'b1, 1'b0};
4938: data_out = {8'd67, 8'd147, 1'b1, 1'b0};
4939: data_out = {8'd77, 8'd147, 1'b1, 1'b0};
4940: data_out = {8'd78, 8'd147, 1'b1, 1'b0};
4941: data_out = {8'd79, 8'd147, 1'b1, 1'b0};
4942: data_out = {8'd80, 8'd147, 1'b1, 1'b0};
4943: data_out = {8'd81, 8'd147, 1'b1, 1'b0};
4944: data_out = {8'd83, 8'd147, 1'b1, 1'b0};
4945: data_out = {8'd88, 8'd147, 1'b1, 1'b0};
4946: data_out = {8'd91, 8'd147, 1'b1, 1'b0};
4947: data_out = {8'd92, 8'd147, 1'b1, 1'b0};
4948: data_out = {8'd93, 8'd147, 1'b1, 1'b0};
4949: data_out = {8'd94, 8'd147, 1'b1, 1'b0};
4950: data_out = {8'd95, 8'd147, 1'b1, 1'b0};
4951: data_out = {8'd100, 8'd147, 1'b1, 1'b0};
4952: data_out = {8'd105, 8'd147, 1'b1, 1'b0};
4953: data_out = {8'd115, 8'd147, 1'b1, 1'b0};
4954: data_out = {8'd116, 8'd147, 1'b1, 1'b0};
4955: data_out = {8'd117, 8'd147, 1'b1, 1'b0};
4956: data_out = {8'd118, 8'd147, 1'b1, 1'b0};
4957: data_out = {8'd119, 8'd147, 1'b1, 1'b0};
4958: data_out = {8'd121, 8'd147, 1'b1, 1'b0};
4959: data_out = {8'd126, 8'd147, 1'b1, 1'b0};
4960: data_out = {8'd129, 8'd147, 1'b1, 1'b0};
4961: data_out = {8'd130, 8'd147, 1'b1, 1'b0};
4962: data_out = {8'd131, 8'd147, 1'b1, 1'b0};
4963: data_out = {8'd132, 8'd147, 1'b1, 1'b0};
4964: data_out = {8'd133, 8'd147, 1'b1, 1'b0};
4965: data_out = {8'd135, 8'd147, 1'b1, 1'b0};
4966: data_out = {8'd136, 8'd147, 1'b1, 1'b0};
4967: data_out = {8'd137, 8'd147, 1'b1, 1'b0};
4968: data_out = {8'd138, 8'd147, 1'b1, 1'b0};
4969: data_out = {8'd143, 8'd147, 1'b1, 1'b0};
4970: data_out = {8'd153, 8'd147, 1'b1, 1'b0};
4971: data_out = {8'd154, 8'd147, 1'b1, 1'b0};
4972: data_out = {8'd155, 8'd147, 1'b1, 1'b0};
4973: data_out = {8'd156, 8'd147, 1'b1, 1'b0};
4974: data_out = {8'd157, 8'd147, 1'b1, 1'b0};
4975: data_out = {8'd159, 8'd147, 1'b1, 1'b0};
4976: data_out = {8'd164, 8'd147, 1'b1, 1'b0};
4977: data_out = {8'd167, 8'd147, 1'b1, 1'b0};
4978: data_out = {8'd168, 8'd147, 1'b1, 1'b0};
4979: data_out = {8'd169, 8'd147, 1'b1, 1'b0};
4980: data_out = {8'd170, 8'd147, 1'b1, 1'b0};
4981: data_out = {8'd171, 8'd147, 1'b1, 1'b0};
4982: data_out = {8'd173, 8'd147, 1'b1, 1'b0};
4983: data_out = {8'd174, 8'd147, 1'b1, 1'b0};
4984: data_out = {8'd175, 8'd147, 1'b1, 1'b0};
4985: data_out = {8'd176, 8'd147, 1'b1, 1'b0};
4986: data_out = {8'd177, 8'd147, 1'b1, 1'b0};
4987: data_out = {8'd186, 8'd147, 1'b1, 1'b0};
4988: data_out = {8'd187, 8'd147, 1'b1, 1'b0};
4989: data_out = {8'd188, 8'd147, 1'b1, 1'b0};
4990: data_out = {8'd189, 8'd147, 1'b1, 1'b0};
4991: data_out = {8'd190, 8'd147, 1'b1, 1'b0};
4992: data_out = {8'd193, 8'd147, 1'b1, 1'b0};
4993: data_out = {8'd194, 8'd147, 1'b1, 1'b0};
4994: data_out = {8'd195, 8'd147, 1'b1, 1'b0};
4995: data_out = {8'd196, 8'd147, 1'b1, 1'b0};
4996: data_out = {8'd197, 8'd147, 1'b1, 1'b0};
4997: data_out = {8'd25, 8'd148, 1'b1, 1'b0};
4998: data_out = {8'd66, 8'd148, 1'b1, 1'b0};
4999: data_out = {8'd67, 8'd148, 1'b1, 1'b0};
5000: data_out = {8'd104, 8'd148, 1'b1, 1'b0};
5001: data_out = {8'd105, 8'd148, 1'b1, 1'b0};
5002: data_out = {8'd142, 8'd148, 1'b1, 1'b0};
5003: data_out = {8'd143, 8'd148, 1'b1, 1'b0};
5004: data_out = {8'd193, 8'd148, 1'b1, 1'b0};
5005: data_out = {8'd25, 8'd149, 1'b1, 1'b0};
5006: data_out = {8'd193, 8'd149, 1'b1, 1'b0};
5007: data_out = {8'd25, 8'd150, 1'b1, 1'b0};
5008: data_out = {8'd193, 8'd150, 1'b1, 1'b0};
5009: data_out = {8'd27, 8'd152, 1'b1, 1'b0};
5010: data_out = {8'd40, 8'd152, 1'b1, 1'b0};
5011: data_out = {8'd52, 8'd152, 1'b1, 1'b0};
5012: data_out = {8'd63, 8'd152, 1'b1, 1'b0};
5013: data_out = {8'd64, 8'd152, 1'b1, 1'b0};
5014: data_out = {8'd65, 8'd152, 1'b1, 1'b0};
5015: data_out = {8'd71, 8'd152, 1'b1, 1'b0};
5016: data_out = {8'd127, 8'd152, 1'b1, 1'b0};
5017: data_out = {8'd6, 8'd153, 1'b1, 1'b0};
5018: data_out = {8'd44, 8'd153, 1'b1, 1'b0};
5019: data_out = {8'd65, 8'd153, 1'b1, 1'b0};
5020: data_out = {8'd127, 8'd153, 1'b1, 1'b0};
5021: data_out = {8'd5, 8'd154, 1'b1, 1'b0};
5022: data_out = {8'd6, 8'd154, 1'b1, 1'b0};
5023: data_out = {8'd7, 8'd154, 1'b1, 1'b0};
5024: data_out = {8'd8, 8'd154, 1'b1, 1'b0};
5025: data_out = {8'd9, 8'd154, 1'b1, 1'b0};
5026: data_out = {8'd12, 8'd154, 1'b1, 1'b0};
5027: data_out = {8'd13, 8'd154, 1'b1, 1'b0};
5028: data_out = {8'd14, 8'd154, 1'b1, 1'b0};
5029: data_out = {8'd15, 8'd154, 1'b1, 1'b0};
5030: data_out = {8'd16, 8'd154, 1'b1, 1'b0};
5031: data_out = {8'd25, 8'd154, 1'b1, 1'b0};
5032: data_out = {8'd26, 8'd154, 1'b1, 1'b0};
5033: data_out = {8'd27, 8'd154, 1'b1, 1'b0};
5034: data_out = {8'd31, 8'd154, 1'b1, 1'b0};
5035: data_out = {8'd32, 8'd154, 1'b1, 1'b0};
5036: data_out = {8'd33, 8'd154, 1'b1, 1'b0};
5037: data_out = {8'd34, 8'd154, 1'b1, 1'b0};
5038: data_out = {8'd35, 8'd154, 1'b1, 1'b0};
5039: data_out = {8'd38, 8'd154, 1'b1, 1'b0};
5040: data_out = {8'd39, 8'd154, 1'b1, 1'b0};
5041: data_out = {8'd40, 8'd154, 1'b1, 1'b0};
5042: data_out = {8'd43, 8'd154, 1'b1, 1'b0};
5043: data_out = {8'd44, 8'd154, 1'b1, 1'b0};
5044: data_out = {8'd45, 8'd154, 1'b1, 1'b0};
5045: data_out = {8'd46, 8'd154, 1'b1, 1'b0};
5046: data_out = {8'd47, 8'd154, 1'b1, 1'b0};
5047: data_out = {8'd50, 8'd154, 1'b1, 1'b0};
5048: data_out = {8'd51, 8'd154, 1'b1, 1'b0};
5049: data_out = {8'd52, 8'd154, 1'b1, 1'b0};
5050: data_out = {8'd56, 8'd154, 1'b1, 1'b0};
5051: data_out = {8'd57, 8'd154, 1'b1, 1'b0};
5052: data_out = {8'd58, 8'd154, 1'b1, 1'b0};
5053: data_out = {8'd59, 8'd154, 1'b1, 1'b0};
5054: data_out = {8'd60, 8'd154, 1'b1, 1'b0};
5055: data_out = {8'd65, 8'd154, 1'b1, 1'b0};
5056: data_out = {8'd69, 8'd154, 1'b1, 1'b0};
5057: data_out = {8'd70, 8'd154, 1'b1, 1'b0};
5058: data_out = {8'd71, 8'd154, 1'b1, 1'b0};
5059: data_out = {8'd75, 8'd154, 1'b1, 1'b0};
5060: data_out = {8'd76, 8'd154, 1'b1, 1'b0};
5061: data_out = {8'd77, 8'd154, 1'b1, 1'b0};
5062: data_out = {8'd78, 8'd154, 1'b1, 1'b0};
5063: data_out = {8'd79, 8'd154, 1'b1, 1'b0};
5064: data_out = {8'd81, 8'd154, 1'b1, 1'b0};
5065: data_out = {8'd82, 8'd154, 1'b1, 1'b0};
5066: data_out = {8'd83, 8'd154, 1'b1, 1'b0};
5067: data_out = {8'd84, 8'd154, 1'b1, 1'b0};
5068: data_out = {8'd85, 8'd154, 1'b1, 1'b0};
5069: data_out = {8'd94, 8'd154, 1'b1, 1'b0};
5070: data_out = {8'd98, 8'd154, 1'b1, 1'b0};
5071: data_out = {8'd101, 8'd154, 1'b1, 1'b0};
5072: data_out = {8'd102, 8'd154, 1'b1, 1'b0};
5073: data_out = {8'd103, 8'd154, 1'b1, 1'b0};
5074: data_out = {8'd104, 8'd154, 1'b1, 1'b0};
5075: data_out = {8'd105, 8'd154, 1'b1, 1'b0};
5076: data_out = {8'd108, 8'd154, 1'b1, 1'b0};
5077: data_out = {8'd112, 8'd154, 1'b1, 1'b0};
5078: data_out = {8'd116, 8'd154, 1'b1, 1'b0};
5079: data_out = {8'd117, 8'd154, 1'b1, 1'b0};
5080: data_out = {8'd118, 8'd154, 1'b1, 1'b0};
5081: data_out = {8'd127, 8'd154, 1'b1, 1'b0};
5082: data_out = {8'd128, 8'd154, 1'b1, 1'b0};
5083: data_out = {8'd129, 8'd154, 1'b1, 1'b0};
5084: data_out = {8'd130, 8'd154, 1'b1, 1'b0};
5085: data_out = {8'd131, 8'd154, 1'b1, 1'b0};
5086: data_out = {8'd134, 8'd154, 1'b1, 1'b0};
5087: data_out = {8'd135, 8'd154, 1'b1, 1'b0};
5088: data_out = {8'd136, 8'd154, 1'b1, 1'b0};
5089: data_out = {8'd137, 8'd154, 1'b1, 1'b0};
5090: data_out = {8'd138, 8'd154, 1'b1, 1'b0};
5091: data_out = {8'd141, 8'd154, 1'b1, 1'b0};
5092: data_out = {8'd142, 8'd154, 1'b1, 1'b0};
5093: data_out = {8'd143, 8'd154, 1'b1, 1'b0};
5094: data_out = {8'd144, 8'd154, 1'b1, 1'b0};
5095: data_out = {8'd145, 8'd154, 1'b1, 1'b0};
5096: data_out = {8'd148, 8'd154, 1'b1, 1'b0};
5097: data_out = {8'd152, 8'd154, 1'b1, 1'b0};
5098: data_out = {8'd155, 8'd154, 1'b1, 1'b0};
5099: data_out = {8'd156, 8'd154, 1'b1, 1'b0};
5100: data_out = {8'd157, 8'd154, 1'b1, 1'b0};
5101: data_out = {8'd158, 8'd154, 1'b1, 1'b0};
5102: data_out = {8'd159, 8'd154, 1'b1, 1'b0};
5103: data_out = {8'd162, 8'd154, 1'b1, 1'b0};
5104: data_out = {8'd163, 8'd154, 1'b1, 1'b0};
5105: data_out = {8'd164, 8'd154, 1'b1, 1'b0};
5106: data_out = {8'd165, 8'd154, 1'b1, 1'b0};
5107: data_out = {8'd6, 8'd155, 1'b1, 1'b0};
5108: data_out = {8'd12, 8'd155, 1'b1, 1'b0};
5109: data_out = {8'd16, 8'd155, 1'b1, 1'b0};
5110: data_out = {8'd27, 8'd155, 1'b1, 1'b0};
5111: data_out = {8'd31, 8'd155, 1'b1, 1'b0};
5112: data_out = {8'd35, 8'd155, 1'b1, 1'b0};
5113: data_out = {8'd40, 8'd155, 1'b1, 1'b0};
5114: data_out = {8'd44, 8'd155, 1'b1, 1'b0};
5115: data_out = {8'd52, 8'd155, 1'b1, 1'b0};
5116: data_out = {8'd56, 8'd155, 1'b1, 1'b0};
5117: data_out = {8'd60, 8'd155, 1'b1, 1'b0};
5118: data_out = {8'd65, 8'd155, 1'b1, 1'b0};
5119: data_out = {8'd71, 8'd155, 1'b1, 1'b0};
5120: data_out = {8'd75, 8'd155, 1'b1, 1'b0};
5121: data_out = {8'd78, 8'd155, 1'b1, 1'b0};
5122: data_out = {8'd81, 8'd155, 1'b1, 1'b0};
5123: data_out = {8'd85, 8'd155, 1'b1, 1'b0};
5124: data_out = {8'd94, 8'd155, 1'b1, 1'b0};
5125: data_out = {8'd98, 8'd155, 1'b1, 1'b0};
5126: data_out = {8'd101, 8'd155, 1'b1, 1'b0};
5127: data_out = {8'd105, 8'd155, 1'b1, 1'b0};
5128: data_out = {8'd108, 8'd155, 1'b1, 1'b0};
5129: data_out = {8'd112, 8'd155, 1'b1, 1'b0};
5130: data_out = {8'd116, 8'd155, 1'b1, 1'b0};
5131: data_out = {8'd118, 8'd155, 1'b1, 1'b0};
5132: data_out = {8'd127, 8'd155, 1'b1, 1'b0};
5133: data_out = {8'd131, 8'd155, 1'b1, 1'b0};
5134: data_out = {8'd134, 8'd155, 1'b1, 1'b0};
5135: data_out = {8'd138, 8'd155, 1'b1, 1'b0};
5136: data_out = {8'd141, 8'd155, 1'b1, 1'b0};
5137: data_out = {8'd145, 8'd155, 1'b1, 1'b0};
5138: data_out = {8'd148, 8'd155, 1'b1, 1'b0};
5139: data_out = {8'd152, 8'd155, 1'b1, 1'b0};
5140: data_out = {8'd155, 8'd155, 1'b1, 1'b0};
5141: data_out = {8'd159, 8'd155, 1'b1, 1'b0};
5142: data_out = {8'd162, 8'd155, 1'b1, 1'b0};
5143: data_out = {8'd165, 8'd155, 1'b1, 1'b0};
5144: data_out = {8'd6, 8'd156, 1'b1, 1'b0};
5145: data_out = {8'd12, 8'd156, 1'b1, 1'b0};
5146: data_out = {8'd16, 8'd156, 1'b1, 1'b0};
5147: data_out = {8'd27, 8'd156, 1'b1, 1'b0};
5148: data_out = {8'd31, 8'd156, 1'b1, 1'b0};
5149: data_out = {8'd35, 8'd156, 1'b1, 1'b0};
5150: data_out = {8'd40, 8'd156, 1'b1, 1'b0};
5151: data_out = {8'd44, 8'd156, 1'b1, 1'b0};
5152: data_out = {8'd52, 8'd156, 1'b1, 1'b0};
5153: data_out = {8'd60, 8'd156, 1'b1, 1'b0};
5154: data_out = {8'd65, 8'd156, 1'b1, 1'b0};
5155: data_out = {8'd71, 8'd156, 1'b1, 1'b0};
5156: data_out = {8'd78, 8'd156, 1'b1, 1'b0};
5157: data_out = {8'd81, 8'd156, 1'b1, 1'b0};
5158: data_out = {8'd85, 8'd156, 1'b1, 1'b0};
5159: data_out = {8'd94, 8'd156, 1'b1, 1'b0};
5160: data_out = {8'd98, 8'd156, 1'b1, 1'b0};
5161: data_out = {8'd101, 8'd156, 1'b1, 1'b0};
5162: data_out = {8'd105, 8'd156, 1'b1, 1'b0};
5163: data_out = {8'd108, 8'd156, 1'b1, 1'b0};
5164: data_out = {8'd112, 8'd156, 1'b1, 1'b0};
5165: data_out = {8'd116, 8'd156, 1'b1, 1'b0};
5166: data_out = {8'd127, 8'd156, 1'b1, 1'b0};
5167: data_out = {8'd131, 8'd156, 1'b1, 1'b0};
5168: data_out = {8'd138, 8'd156, 1'b1, 1'b0};
5169: data_out = {8'd141, 8'd156, 1'b1, 1'b0};
5170: data_out = {8'd148, 8'd156, 1'b1, 1'b0};
5171: data_out = {8'd152, 8'd156, 1'b1, 1'b0};
5172: data_out = {8'd155, 8'd156, 1'b1, 1'b0};
5173: data_out = {8'd164, 8'd156, 1'b1, 1'b0};
5174: data_out = {8'd6, 8'd157, 1'b1, 1'b0};
5175: data_out = {8'd12, 8'd157, 1'b1, 1'b0};
5176: data_out = {8'd16, 8'd157, 1'b1, 1'b0};
5177: data_out = {8'd27, 8'd157, 1'b1, 1'b0};
5178: data_out = {8'd31, 8'd157, 1'b1, 1'b0};
5179: data_out = {8'd35, 8'd157, 1'b1, 1'b0};
5180: data_out = {8'd40, 8'd157, 1'b1, 1'b0};
5181: data_out = {8'd44, 8'd157, 1'b1, 1'b0};
5182: data_out = {8'd52, 8'd157, 1'b1, 1'b0};
5183: data_out = {8'd57, 8'd157, 1'b1, 1'b0};
5184: data_out = {8'd58, 8'd157, 1'b1, 1'b0};
5185: data_out = {8'd59, 8'd157, 1'b1, 1'b0};
5186: data_out = {8'd60, 8'd157, 1'b1, 1'b0};
5187: data_out = {8'd65, 8'd157, 1'b1, 1'b0};
5188: data_out = {8'd71, 8'd157, 1'b1, 1'b0};
5189: data_out = {8'd77, 8'd157, 1'b1, 1'b0};
5190: data_out = {8'd81, 8'd157, 1'b1, 1'b0};
5191: data_out = {8'd82, 8'd157, 1'b1, 1'b0};
5192: data_out = {8'd83, 8'd157, 1'b1, 1'b0};
5193: data_out = {8'd84, 8'd157, 1'b1, 1'b0};
5194: data_out = {8'd94, 8'd157, 1'b1, 1'b0};
5195: data_out = {8'd98, 8'd157, 1'b1, 1'b0};
5196: data_out = {8'd101, 8'd157, 1'b1, 1'b0};
5197: data_out = {8'd105, 8'd157, 1'b1, 1'b0};
5198: data_out = {8'd108, 8'd157, 1'b1, 1'b0};
5199: data_out = {8'd112, 8'd157, 1'b1, 1'b0};
5200: data_out = {8'd116, 8'd157, 1'b1, 1'b0};
5201: data_out = {8'd127, 8'd157, 1'b1, 1'b0};
5202: data_out = {8'd131, 8'd157, 1'b1, 1'b0};
5203: data_out = {8'd135, 8'd157, 1'b1, 1'b0};
5204: data_out = {8'd136, 8'd157, 1'b1, 1'b0};
5205: data_out = {8'd137, 8'd157, 1'b1, 1'b0};
5206: data_out = {8'd138, 8'd157, 1'b1, 1'b0};
5207: data_out = {8'd141, 8'd157, 1'b1, 1'b0};
5208: data_out = {8'd142, 8'd157, 1'b1, 1'b0};
5209: data_out = {8'd143, 8'd157, 1'b1, 1'b0};
5210: data_out = {8'd144, 8'd157, 1'b1, 1'b0};
5211: data_out = {8'd145, 8'd157, 1'b1, 1'b0};
5212: data_out = {8'd148, 8'd157, 1'b1, 1'b0};
5213: data_out = {8'd152, 8'd157, 1'b1, 1'b0};
5214: data_out = {8'd155, 8'd157, 1'b1, 1'b0};
5215: data_out = {8'd156, 8'd157, 1'b1, 1'b0};
5216: data_out = {8'd157, 8'd157, 1'b1, 1'b0};
5217: data_out = {8'd158, 8'd157, 1'b1, 1'b0};
5218: data_out = {8'd159, 8'd157, 1'b1, 1'b0};
5219: data_out = {8'd163, 8'd157, 1'b1, 1'b0};
5220: data_out = {8'd164, 8'd157, 1'b1, 1'b0};
5221: data_out = {8'd165, 8'd157, 1'b1, 1'b0};
5222: data_out = {8'd6, 8'd158, 1'b1, 1'b0};
5223: data_out = {8'd12, 8'd158, 1'b1, 1'b0};
5224: data_out = {8'd16, 8'd158, 1'b1, 1'b0};
5225: data_out = {8'd27, 8'd158, 1'b1, 1'b0};
5226: data_out = {8'd31, 8'd158, 1'b1, 1'b0};
5227: data_out = {8'd35, 8'd158, 1'b1, 1'b0};
5228: data_out = {8'd40, 8'd158, 1'b1, 1'b0};
5229: data_out = {8'd44, 8'd158, 1'b1, 1'b0};
5230: data_out = {8'd52, 8'd158, 1'b1, 1'b0};
5231: data_out = {8'd56, 8'd158, 1'b1, 1'b0};
5232: data_out = {8'd60, 8'd158, 1'b1, 1'b0};
5233: data_out = {8'd65, 8'd158, 1'b1, 1'b0};
5234: data_out = {8'd71, 8'd158, 1'b1, 1'b0};
5235: data_out = {8'd76, 8'd158, 1'b1, 1'b0};
5236: data_out = {8'd81, 8'd158, 1'b1, 1'b0};
5237: data_out = {8'd94, 8'd158, 1'b1, 1'b0};
5238: data_out = {8'd98, 8'd158, 1'b1, 1'b0};
5239: data_out = {8'd101, 8'd158, 1'b1, 1'b0};
5240: data_out = {8'd105, 8'd158, 1'b1, 1'b0};
5241: data_out = {8'd108, 8'd158, 1'b1, 1'b0};
5242: data_out = {8'd112, 8'd158, 1'b1, 1'b0};
5243: data_out = {8'd116, 8'd158, 1'b1, 1'b0};
5244: data_out = {8'd127, 8'd158, 1'b1, 1'b0};
5245: data_out = {8'd131, 8'd158, 1'b1, 1'b0};
5246: data_out = {8'd134, 8'd158, 1'b1, 1'b0};
5247: data_out = {8'd138, 8'd158, 1'b1, 1'b0};
5248: data_out = {8'd145, 8'd158, 1'b1, 1'b0};
5249: data_out = {8'd148, 8'd158, 1'b1, 1'b0};
5250: data_out = {8'd152, 8'd158, 1'b1, 1'b0};
5251: data_out = {8'd159, 8'd158, 1'b1, 1'b0};
5252: data_out = {8'd165, 8'd158, 1'b1, 1'b0};
5253: data_out = {8'd6, 8'd159, 1'b1, 1'b0};
5254: data_out = {8'd12, 8'd159, 1'b1, 1'b0};
5255: data_out = {8'd16, 8'd159, 1'b1, 1'b0};
5256: data_out = {8'd27, 8'd159, 1'b1, 1'b0};
5257: data_out = {8'd31, 8'd159, 1'b1, 1'b0};
5258: data_out = {8'd35, 8'd159, 1'b1, 1'b0};
5259: data_out = {8'd40, 8'd159, 1'b1, 1'b0};
5260: data_out = {8'd44, 8'd159, 1'b1, 1'b0};
5261: data_out = {8'd52, 8'd159, 1'b1, 1'b0};
5262: data_out = {8'd56, 8'd159, 1'b1, 1'b0};
5263: data_out = {8'd60, 8'd159, 1'b1, 1'b0};
5264: data_out = {8'd65, 8'd159, 1'b1, 1'b0};
5265: data_out = {8'd71, 8'd159, 1'b1, 1'b0};
5266: data_out = {8'd75, 8'd159, 1'b1, 1'b0};
5267: data_out = {8'd81, 8'd159, 1'b1, 1'b0};
5268: data_out = {8'd94, 8'd159, 1'b1, 1'b0};
5269: data_out = {8'd98, 8'd159, 1'b1, 1'b0};
5270: data_out = {8'd101, 8'd159, 1'b1, 1'b0};
5271: data_out = {8'd105, 8'd159, 1'b1, 1'b0};
5272: data_out = {8'd108, 8'd159, 1'b1, 1'b0};
5273: data_out = {8'd112, 8'd159, 1'b1, 1'b0};
5274: data_out = {8'd116, 8'd159, 1'b1, 1'b0};
5275: data_out = {8'd127, 8'd159, 1'b1, 1'b0};
5276: data_out = {8'd131, 8'd159, 1'b1, 1'b0};
5277: data_out = {8'd134, 8'd159, 1'b1, 1'b0};
5278: data_out = {8'd138, 8'd159, 1'b1, 1'b0};
5279: data_out = {8'd145, 8'd159, 1'b1, 1'b0};
5280: data_out = {8'd148, 8'd159, 1'b1, 1'b0};
5281: data_out = {8'd152, 8'd159, 1'b1, 1'b0};
5282: data_out = {8'd159, 8'd159, 1'b1, 1'b0};
5283: data_out = {8'd165, 8'd159, 1'b1, 1'b0};
5284: data_out = {8'd6, 8'd160, 1'b1, 1'b0};
5285: data_out = {8'd7, 8'd160, 1'b1, 1'b0};
5286: data_out = {8'd8, 8'd160, 1'b1, 1'b0};
5287: data_out = {8'd9, 8'd160, 1'b1, 1'b0};
5288: data_out = {8'd10, 8'd160, 1'b1, 1'b0};
5289: data_out = {8'd12, 8'd160, 1'b1, 1'b0};
5290: data_out = {8'd13, 8'd160, 1'b1, 1'b0};
5291: data_out = {8'd14, 8'd160, 1'b1, 1'b0};
5292: data_out = {8'd15, 8'd160, 1'b1, 1'b0};
5293: data_out = {8'd16, 8'd160, 1'b1, 1'b0};
5294: data_out = {8'd25, 8'd160, 1'b1, 1'b0};
5295: data_out = {8'd26, 8'd160, 1'b1, 1'b0};
5296: data_out = {8'd27, 8'd160, 1'b1, 1'b0};
5297: data_out = {8'd28, 8'd160, 1'b1, 1'b0};
5298: data_out = {8'd29, 8'd160, 1'b1, 1'b0};
5299: data_out = {8'd31, 8'd160, 1'b1, 1'b0};
5300: data_out = {8'd35, 8'd160, 1'b1, 1'b0};
5301: data_out = {8'd38, 8'd160, 1'b1, 1'b0};
5302: data_out = {8'd39, 8'd160, 1'b1, 1'b0};
5303: data_out = {8'd40, 8'd160, 1'b1, 1'b0};
5304: data_out = {8'd41, 8'd160, 1'b1, 1'b0};
5305: data_out = {8'd42, 8'd160, 1'b1, 1'b0};
5306: data_out = {8'd44, 8'd160, 1'b1, 1'b0};
5307: data_out = {8'd45, 8'd160, 1'b1, 1'b0};
5308: data_out = {8'd46, 8'd160, 1'b1, 1'b0};
5309: data_out = {8'd47, 8'd160, 1'b1, 1'b0};
5310: data_out = {8'd48, 8'd160, 1'b1, 1'b0};
5311: data_out = {8'd50, 8'd160, 1'b1, 1'b0};
5312: data_out = {8'd51, 8'd160, 1'b1, 1'b0};
5313: data_out = {8'd52, 8'd160, 1'b1, 1'b0};
5314: data_out = {8'd53, 8'd160, 1'b1, 1'b0};
5315: data_out = {8'd54, 8'd160, 1'b1, 1'b0};
5316: data_out = {8'd56, 8'd160, 1'b1, 1'b0};
5317: data_out = {8'd57, 8'd160, 1'b1, 1'b0};
5318: data_out = {8'd58, 8'd160, 1'b1, 1'b0};
5319: data_out = {8'd59, 8'd160, 1'b1, 1'b0};
5320: data_out = {8'd60, 8'd160, 1'b1, 1'b0};
5321: data_out = {8'd63, 8'd160, 1'b1, 1'b0};
5322: data_out = {8'd64, 8'd160, 1'b1, 1'b0};
5323: data_out = {8'd65, 8'd160, 1'b1, 1'b0};
5324: data_out = {8'd66, 8'd160, 1'b1, 1'b0};
5325: data_out = {8'd67, 8'd160, 1'b1, 1'b0};
5326: data_out = {8'd69, 8'd160, 1'b1, 1'b0};
5327: data_out = {8'd70, 8'd160, 1'b1, 1'b0};
5328: data_out = {8'd71, 8'd160, 1'b1, 1'b0};
5329: data_out = {8'd72, 8'd160, 1'b1, 1'b0};
5330: data_out = {8'd73, 8'd160, 1'b1, 1'b0};
5331: data_out = {8'd75, 8'd160, 1'b1, 1'b0};
5332: data_out = {8'd76, 8'd160, 1'b1, 1'b0};
5333: data_out = {8'd77, 8'd160, 1'b1, 1'b0};
5334: data_out = {8'd78, 8'd160, 1'b1, 1'b0};
5335: data_out = {8'd79, 8'd160, 1'b1, 1'b0};
5336: data_out = {8'd81, 8'd160, 1'b1, 1'b0};
5337: data_out = {8'd82, 8'd160, 1'b1, 1'b0};
5338: data_out = {8'd83, 8'd160, 1'b1, 1'b0};
5339: data_out = {8'd84, 8'd160, 1'b1, 1'b0};
5340: data_out = {8'd85, 8'd160, 1'b1, 1'b0};
5341: data_out = {8'd94, 8'd160, 1'b1, 1'b0};
5342: data_out = {8'd95, 8'd160, 1'b1, 1'b0};
5343: data_out = {8'd96, 8'd160, 1'b1, 1'b0};
5344: data_out = {8'd97, 8'd160, 1'b1, 1'b0};
5345: data_out = {8'd98, 8'd160, 1'b1, 1'b0};
5346: data_out = {8'd101, 8'd160, 1'b1, 1'b0};
5347: data_out = {8'd102, 8'd160, 1'b1, 1'b0};
5348: data_out = {8'd103, 8'd160, 1'b1, 1'b0};
5349: data_out = {8'd104, 8'd160, 1'b1, 1'b0};
5350: data_out = {8'd105, 8'd160, 1'b1, 1'b0};
5351: data_out = {8'd108, 8'd160, 1'b1, 1'b0};
5352: data_out = {8'd109, 8'd160, 1'b1, 1'b0};
5353: data_out = {8'd110, 8'd160, 1'b1, 1'b0};
5354: data_out = {8'd111, 8'd160, 1'b1, 1'b0};
5355: data_out = {8'd112, 8'd160, 1'b1, 1'b0};
5356: data_out = {8'd114, 8'd160, 1'b1, 1'b0};
5357: data_out = {8'd115, 8'd160, 1'b1, 1'b0};
5358: data_out = {8'd116, 8'd160, 1'b1, 1'b0};
5359: data_out = {8'd117, 8'd160, 1'b1, 1'b0};
5360: data_out = {8'd118, 8'd160, 1'b1, 1'b0};
5361: data_out = {8'd119, 8'd160, 1'b1, 1'b0};
5362: data_out = {8'd127, 8'd160, 1'b1, 1'b0};
5363: data_out = {8'd128, 8'd160, 1'b1, 1'b0};
5364: data_out = {8'd129, 8'd160, 1'b1, 1'b0};
5365: data_out = {8'd130, 8'd160, 1'b1, 1'b0};
5366: data_out = {8'd131, 8'd160, 1'b1, 1'b0};
5367: data_out = {8'd134, 8'd160, 1'b1, 1'b0};
5368: data_out = {8'd135, 8'd160, 1'b1, 1'b0};
5369: data_out = {8'd136, 8'd160, 1'b1, 1'b0};
5370: data_out = {8'd137, 8'd160, 1'b1, 1'b0};
5371: data_out = {8'd138, 8'd160, 1'b1, 1'b0};
5372: data_out = {8'd141, 8'd160, 1'b1, 1'b0};
5373: data_out = {8'd142, 8'd160, 1'b1, 1'b0};
5374: data_out = {8'd143, 8'd160, 1'b1, 1'b0};
5375: data_out = {8'd144, 8'd160, 1'b1, 1'b0};
5376: data_out = {8'd145, 8'd160, 1'b1, 1'b0};
5377: data_out = {8'd148, 8'd160, 1'b1, 1'b0};
5378: data_out = {8'd149, 8'd160, 1'b1, 1'b0};
5379: data_out = {8'd150, 8'd160, 1'b1, 1'b0};
5380: data_out = {8'd151, 8'd160, 1'b1, 1'b0};
5381: data_out = {8'd152, 8'd160, 1'b1, 1'b0};
5382: data_out = {8'd155, 8'd160, 1'b1, 1'b0};
5383: data_out = {8'd156, 8'd160, 1'b1, 1'b0};
5384: data_out = {8'd157, 8'd160, 1'b1, 1'b0};
5385: data_out = {8'd158, 8'd160, 1'b1, 1'b0};
5386: data_out = {8'd159, 8'd160, 1'b1, 1'b0};
5387: data_out = {8'd162, 8'd160, 1'b1, 1'b0};
5388: data_out = {8'd163, 8'd160, 1'b1, 1'b0};
5389: data_out = {8'd164, 8'd160, 1'b1, 1'b0};
5390: data_out = {8'd165, 8'd160, 1'b1, 1'b0};
5391: data_out = {8'd98, 8'd161, 1'b1, 1'b0};
5392: data_out = {8'd152, 8'd161, 1'b1, 1'b0};
5393: data_out = {8'd98, 8'd162, 1'b1, 1'b0};
5394: data_out = {8'd152, 8'd162, 1'b1, 1'b0};
5395: data_out = {8'd94, 8'd163, 1'b1, 1'b0};
5396: data_out = {8'd95, 8'd163, 1'b1, 1'b0};
5397: data_out = {8'd96, 8'd163, 1'b1, 1'b0};
5398: data_out = {8'd97, 8'd163, 1'b1, 1'b0};
5399: data_out = {8'd98, 8'd163, 1'b1, 1'b0};
5400: data_out = {8'd148, 8'd163, 1'b1, 1'b0};
5401: data_out = {8'd149, 8'd163, 1'b1, 1'b0};
5402: data_out = {8'd150, 8'd163, 1'b1, 1'b0};
5403: data_out = {8'd151, 8'd163, 1'b1, 1'b0};
5404: data_out = {8'd152, 8'd163, 1'b1, 1'b0};
5405: data_out = {8'd101, 8'd164, 1'b1, 1'b0};
5406: data_out = {8'd102, 8'd164, 1'b1, 1'b0};
5407: data_out = {8'd103, 8'd164, 1'b1, 1'b0};
5408: data_out = {8'd104, 8'd164, 1'b1, 1'b0};
5409: data_out = {8'd70, 8'd165, 1'b1, 1'b0};
5410: data_out = {8'd90, 8'd165, 1'b1, 1'b0};
5411: data_out = {8'd101, 8'd165, 1'b1, 1'b0};
5412: data_out = {8'd104, 8'd165, 1'b1, 1'b0};
5413: data_out = {8'd49, 8'd166, 1'b1, 1'b0};
5414: data_out = {8'd90, 8'd166, 1'b1, 1'b0};
5415: data_out = {8'd101, 8'd166, 1'b1, 1'b0};
5416: data_out = {8'd162, 8'd166, 1'b1, 1'b0};
5417: data_out = {8'd6, 8'd167, 1'b1, 1'b0};
5418: data_out = {8'd7, 8'd167, 1'b1, 1'b0};
5419: data_out = {8'd8, 8'd167, 1'b1, 1'b0};
5420: data_out = {8'd9, 8'd167, 1'b1, 1'b0};
5421: data_out = {8'd10, 8'd167, 1'b1, 1'b0};
5422: data_out = {8'd13, 8'd167, 1'b1, 1'b0};
5423: data_out = {8'd14, 8'd167, 1'b1, 1'b0};
5424: data_out = {8'd15, 8'd167, 1'b1, 1'b0};
5425: data_out = {8'd16, 8'd167, 1'b1, 1'b0};
5426: data_out = {8'd17, 8'd167, 1'b1, 1'b0};
5427: data_out = {8'd19, 8'd167, 1'b1, 1'b0};
5428: data_out = {8'd20, 8'd167, 1'b1, 1'b0};
5429: data_out = {8'd21, 8'd167, 1'b1, 1'b0};
5430: data_out = {8'd22, 8'd167, 1'b1, 1'b0};
5431: data_out = {8'd23, 8'd167, 1'b1, 1'b0};
5432: data_out = {8'd24, 8'd167, 1'b1, 1'b0};
5433: data_out = {8'd25, 8'd167, 1'b1, 1'b0};
5434: data_out = {8'd28, 8'd167, 1'b1, 1'b0};
5435: data_out = {8'd29, 8'd167, 1'b1, 1'b0};
5436: data_out = {8'd30, 8'd167, 1'b1, 1'b0};
5437: data_out = {8'd31, 8'd167, 1'b1, 1'b0};
5438: data_out = {8'd32, 8'd167, 1'b1, 1'b0};
5439: data_out = {8'd35, 8'd167, 1'b1, 1'b0};
5440: data_out = {8'd36, 8'd167, 1'b1, 1'b0};
5441: data_out = {8'd37, 8'd167, 1'b1, 1'b0};
5442: data_out = {8'd38, 8'd167, 1'b1, 1'b0};
5443: data_out = {8'd39, 8'd167, 1'b1, 1'b0};
5444: data_out = {8'd42, 8'd167, 1'b1, 1'b0};
5445: data_out = {8'd43, 8'd167, 1'b1, 1'b0};
5446: data_out = {8'd44, 8'd167, 1'b1, 1'b0};
5447: data_out = {8'd45, 8'd167, 1'b1, 1'b0};
5448: data_out = {8'd46, 8'd167, 1'b1, 1'b0};
5449: data_out = {8'd48, 8'd167, 1'b1, 1'b0};
5450: data_out = {8'd49, 8'd167, 1'b1, 1'b0};
5451: data_out = {8'd50, 8'd167, 1'b1, 1'b0};
5452: data_out = {8'd51, 8'd167, 1'b1, 1'b0};
5453: data_out = {8'd52, 8'd167, 1'b1, 1'b0};
5454: data_out = {8'd61, 8'd167, 1'b1, 1'b0};
5455: data_out = {8'd62, 8'd167, 1'b1, 1'b0};
5456: data_out = {8'd63, 8'd167, 1'b1, 1'b0};
5457: data_out = {8'd64, 8'd167, 1'b1, 1'b0};
5458: data_out = {8'd65, 8'd167, 1'b1, 1'b0};
5459: data_out = {8'd68, 8'd167, 1'b1, 1'b0};
5460: data_out = {8'd69, 8'd167, 1'b1, 1'b0};
5461: data_out = {8'd70, 8'd167, 1'b1, 1'b0};
5462: data_out = {8'd75, 8'd167, 1'b1, 1'b0};
5463: data_out = {8'd76, 8'd167, 1'b1, 1'b0};
5464: data_out = {8'd77, 8'd167, 1'b1, 1'b0};
5465: data_out = {8'd86, 8'd167, 1'b1, 1'b0};
5466: data_out = {8'd87, 8'd167, 1'b1, 1'b0};
5467: data_out = {8'd88, 8'd167, 1'b1, 1'b0};
5468: data_out = {8'd89, 8'd167, 1'b1, 1'b0};
5469: data_out = {8'd90, 8'd167, 1'b1, 1'b0};
5470: data_out = {8'd93, 8'd167, 1'b1, 1'b0};
5471: data_out = {8'd94, 8'd167, 1'b1, 1'b0};
5472: data_out = {8'd95, 8'd167, 1'b1, 1'b0};
5473: data_out = {8'd96, 8'd167, 1'b1, 1'b0};
5474: data_out = {8'd97, 8'd167, 1'b1, 1'b0};
5475: data_out = {8'd99, 8'd167, 1'b1, 1'b0};
5476: data_out = {8'd100, 8'd167, 1'b1, 1'b0};
5477: data_out = {8'd101, 8'd167, 1'b1, 1'b0};
5478: data_out = {8'd102, 8'd167, 1'b1, 1'b0};
5479: data_out = {8'd103, 8'd167, 1'b1, 1'b0};
5480: data_out = {8'd104, 8'd167, 1'b1, 1'b0};
5481: data_out = {8'd107, 8'd167, 1'b1, 1'b0};
5482: data_out = {8'd108, 8'd167, 1'b1, 1'b0};
5483: data_out = {8'd109, 8'd167, 1'b1, 1'b0};
5484: data_out = {8'd110, 8'd167, 1'b1, 1'b0};
5485: data_out = {8'd111, 8'd167, 1'b1, 1'b0};
5486: data_out = {8'd114, 8'd167, 1'b1, 1'b0};
5487: data_out = {8'd115, 8'd167, 1'b1, 1'b0};
5488: data_out = {8'd116, 8'd167, 1'b1, 1'b0};
5489: data_out = {8'd117, 8'd167, 1'b1, 1'b0};
5490: data_out = {8'd118, 8'd167, 1'b1, 1'b0};
5491: data_out = {8'd121, 8'd167, 1'b1, 1'b0};
5492: data_out = {8'd122, 8'd167, 1'b1, 1'b0};
5493: data_out = {8'd123, 8'd167, 1'b1, 1'b0};
5494: data_out = {8'd124, 8'd167, 1'b1, 1'b0};
5495: data_out = {8'd125, 8'd167, 1'b1, 1'b0};
5496: data_out = {8'd128, 8'd167, 1'b1, 1'b0};
5497: data_out = {8'd129, 8'd167, 1'b1, 1'b0};
5498: data_out = {8'd130, 8'd167, 1'b1, 1'b0};
5499: data_out = {8'd131, 8'd167, 1'b1, 1'b0};
5500: data_out = {8'd132, 8'd167, 1'b1, 1'b0};
5501: data_out = {8'd141, 8'd167, 1'b1, 1'b0};
5502: data_out = {8'd142, 8'd167, 1'b1, 1'b0};
5503: data_out = {8'd143, 8'd167, 1'b1, 1'b0};
5504: data_out = {8'd144, 8'd167, 1'b1, 1'b0};
5505: data_out = {8'd145, 8'd167, 1'b1, 1'b0};
5506: data_out = {8'd148, 8'd167, 1'b1, 1'b0};
5507: data_out = {8'd152, 8'd167, 1'b1, 1'b0};
5508: data_out = {8'd155, 8'd167, 1'b1, 1'b0};
5509: data_out = {8'd156, 8'd167, 1'b1, 1'b0};
5510: data_out = {8'd157, 8'd167, 1'b1, 1'b0};
5511: data_out = {8'd158, 8'd167, 1'b1, 1'b0};
5512: data_out = {8'd159, 8'd167, 1'b1, 1'b0};
5513: data_out = {8'd161, 8'd167, 1'b1, 1'b0};
5514: data_out = {8'd162, 8'd167, 1'b1, 1'b0};
5515: data_out = {8'd163, 8'd167, 1'b1, 1'b0};
5516: data_out = {8'd164, 8'd167, 1'b1, 1'b0};
5517: data_out = {8'd165, 8'd167, 1'b1, 1'b0};
5518: data_out = {8'd168, 8'd167, 1'b1, 1'b0};
5519: data_out = {8'd169, 8'd167, 1'b1, 1'b0};
5520: data_out = {8'd170, 8'd167, 1'b1, 1'b0};
5521: data_out = {8'd171, 8'd167, 1'b1, 1'b0};
5522: data_out = {8'd172, 8'd167, 1'b1, 1'b0};
5523: data_out = {8'd174, 8'd167, 1'b1, 1'b0};
5524: data_out = {8'd175, 8'd167, 1'b1, 1'b0};
5525: data_out = {8'd176, 8'd167, 1'b1, 1'b0};
5526: data_out = {8'd177, 8'd167, 1'b1, 1'b0};
5527: data_out = {8'd178, 8'd167, 1'b1, 1'b0};
5528: data_out = {8'd179, 8'd167, 1'b1, 1'b0};
5529: data_out = {8'd180, 8'd167, 1'b1, 1'b0};
5530: data_out = {8'd6, 8'd168, 1'b1, 1'b0};
5531: data_out = {8'd10, 8'd168, 1'b1, 1'b0};
5532: data_out = {8'd13, 8'd168, 1'b1, 1'b0};
5533: data_out = {8'd17, 8'd168, 1'b1, 1'b0};
5534: data_out = {8'd19, 8'd168, 1'b1, 1'b0};
5535: data_out = {8'd22, 8'd168, 1'b1, 1'b0};
5536: data_out = {8'd25, 8'd168, 1'b1, 1'b0};
5537: data_out = {8'd28, 8'd168, 1'b1, 1'b0};
5538: data_out = {8'd32, 8'd168, 1'b1, 1'b0};
5539: data_out = {8'd35, 8'd168, 1'b1, 1'b0};
5540: data_out = {8'd39, 8'd168, 1'b1, 1'b0};
5541: data_out = {8'd42, 8'd168, 1'b1, 1'b0};
5542: data_out = {8'd46, 8'd168, 1'b1, 1'b0};
5543: data_out = {8'd49, 8'd168, 1'b1, 1'b0};
5544: data_out = {8'd61, 8'd168, 1'b1, 1'b0};
5545: data_out = {8'd65, 8'd168, 1'b1, 1'b0};
5546: data_out = {8'd70, 8'd168, 1'b1, 1'b0};
5547: data_out = {8'd75, 8'd168, 1'b1, 1'b0};
5548: data_out = {8'd77, 8'd168, 1'b1, 1'b0};
5549: data_out = {8'd86, 8'd168, 1'b1, 1'b0};
5550: data_out = {8'd90, 8'd168, 1'b1, 1'b0};
5551: data_out = {8'd93, 8'd168, 1'b1, 1'b0};
5552: data_out = {8'd97, 8'd168, 1'b1, 1'b0};
5553: data_out = {8'd101, 8'd168, 1'b1, 1'b0};
5554: data_out = {8'd107, 8'd168, 1'b1, 1'b0};
5555: data_out = {8'd111, 8'd168, 1'b1, 1'b0};
5556: data_out = {8'd114, 8'd168, 1'b1, 1'b0};
5557: data_out = {8'd118, 8'd168, 1'b1, 1'b0};
5558: data_out = {8'd121, 8'd168, 1'b1, 1'b0};
5559: data_out = {8'd125, 8'd168, 1'b1, 1'b0};
5560: data_out = {8'd128, 8'd168, 1'b1, 1'b0};
5561: data_out = {8'd132, 8'd168, 1'b1, 1'b0};
5562: data_out = {8'd141, 8'd168, 1'b1, 1'b0};
5563: data_out = {8'd145, 8'd168, 1'b1, 1'b0};
5564: data_out = {8'd148, 8'd168, 1'b1, 1'b0};
5565: data_out = {8'd152, 8'd168, 1'b1, 1'b0};
5566: data_out = {8'd155, 8'd168, 1'b1, 1'b0};
5567: data_out = {8'd159, 8'd168, 1'b1, 1'b0};
5568: data_out = {8'd162, 8'd168, 1'b1, 1'b0};
5569: data_out = {8'd168, 8'd168, 1'b1, 1'b0};
5570: data_out = {8'd172, 8'd168, 1'b1, 1'b0};
5571: data_out = {8'd174, 8'd168, 1'b1, 1'b0};
5572: data_out = {8'd177, 8'd168, 1'b1, 1'b0};
5573: data_out = {8'd180, 8'd168, 1'b1, 1'b0};
5574: data_out = {8'd6, 8'd169, 1'b1, 1'b0};
5575: data_out = {8'd13, 8'd169, 1'b1, 1'b0};
5576: data_out = {8'd17, 8'd169, 1'b1, 1'b0};
5577: data_out = {8'd19, 8'd169, 1'b1, 1'b0};
5578: data_out = {8'd22, 8'd169, 1'b1, 1'b0};
5579: data_out = {8'd25, 8'd169, 1'b1, 1'b0};
5580: data_out = {8'd28, 8'd169, 1'b1, 1'b0};
5581: data_out = {8'd32, 8'd169, 1'b1, 1'b0};
5582: data_out = {8'd39, 8'd169, 1'b1, 1'b0};
5583: data_out = {8'd42, 8'd169, 1'b1, 1'b0};
5584: data_out = {8'd49, 8'd169, 1'b1, 1'b0};
5585: data_out = {8'd65, 8'd169, 1'b1, 1'b0};
5586: data_out = {8'd70, 8'd169, 1'b1, 1'b0};
5587: data_out = {8'd75, 8'd169, 1'b1, 1'b0};
5588: data_out = {8'd86, 8'd169, 1'b1, 1'b0};
5589: data_out = {8'd90, 8'd169, 1'b1, 1'b0};
5590: data_out = {8'd93, 8'd169, 1'b1, 1'b0};
5591: data_out = {8'd97, 8'd169, 1'b1, 1'b0};
5592: data_out = {8'd101, 8'd169, 1'b1, 1'b0};
5593: data_out = {8'd107, 8'd169, 1'b1, 1'b0};
5594: data_out = {8'd111, 8'd169, 1'b1, 1'b0};
5595: data_out = {8'd114, 8'd169, 1'b1, 1'b0};
5596: data_out = {8'd118, 8'd169, 1'b1, 1'b0};
5597: data_out = {8'd121, 8'd169, 1'b1, 1'b0};
5598: data_out = {8'd128, 8'd169, 1'b1, 1'b0};
5599: data_out = {8'd132, 8'd169, 1'b1, 1'b0};
5600: data_out = {8'd141, 8'd169, 1'b1, 1'b0};
5601: data_out = {8'd148, 8'd169, 1'b1, 1'b0};
5602: data_out = {8'd152, 8'd169, 1'b1, 1'b0};
5603: data_out = {8'd155, 8'd169, 1'b1, 1'b0};
5604: data_out = {8'd162, 8'd169, 1'b1, 1'b0};
5605: data_out = {8'd168, 8'd169, 1'b1, 1'b0};
5606: data_out = {8'd172, 8'd169, 1'b1, 1'b0};
5607: data_out = {8'd174, 8'd169, 1'b1, 1'b0};
5608: data_out = {8'd177, 8'd169, 1'b1, 1'b0};
5609: data_out = {8'd180, 8'd169, 1'b1, 1'b0};
5610: data_out = {8'd6, 8'd170, 1'b1, 1'b0};
5611: data_out = {8'd13, 8'd170, 1'b1, 1'b0};
5612: data_out = {8'd17, 8'd170, 1'b1, 1'b0};
5613: data_out = {8'd19, 8'd170, 1'b1, 1'b0};
5614: data_out = {8'd22, 8'd170, 1'b1, 1'b0};
5615: data_out = {8'd25, 8'd170, 1'b1, 1'b0};
5616: data_out = {8'd28, 8'd170, 1'b1, 1'b0};
5617: data_out = {8'd32, 8'd170, 1'b1, 1'b0};
5618: data_out = {8'd36, 8'd170, 1'b1, 1'b0};
5619: data_out = {8'd37, 8'd170, 1'b1, 1'b0};
5620: data_out = {8'd38, 8'd170, 1'b1, 1'b0};
5621: data_out = {8'd39, 8'd170, 1'b1, 1'b0};
5622: data_out = {8'd42, 8'd170, 1'b1, 1'b0};
5623: data_out = {8'd49, 8'd170, 1'b1, 1'b0};
5624: data_out = {8'd62, 8'd170, 1'b1, 1'b0};
5625: data_out = {8'd63, 8'd170, 1'b1, 1'b0};
5626: data_out = {8'd64, 8'd170, 1'b1, 1'b0};
5627: data_out = {8'd65, 8'd170, 1'b1, 1'b0};
5628: data_out = {8'd70, 8'd170, 1'b1, 1'b0};
5629: data_out = {8'd75, 8'd170, 1'b1, 1'b0};
5630: data_out = {8'd86, 8'd170, 1'b1, 1'b0};
5631: data_out = {8'd90, 8'd170, 1'b1, 1'b0};
5632: data_out = {8'd93, 8'd170, 1'b1, 1'b0};
5633: data_out = {8'd94, 8'd170, 1'b1, 1'b0};
5634: data_out = {8'd95, 8'd170, 1'b1, 1'b0};
5635: data_out = {8'd96, 8'd170, 1'b1, 1'b0};
5636: data_out = {8'd101, 8'd170, 1'b1, 1'b0};
5637: data_out = {8'd107, 8'd170, 1'b1, 1'b0};
5638: data_out = {8'd108, 8'd170, 1'b1, 1'b0};
5639: data_out = {8'd109, 8'd170, 1'b1, 1'b0};
5640: data_out = {8'd110, 8'd170, 1'b1, 1'b0};
5641: data_out = {8'd114, 8'd170, 1'b1, 1'b0};
5642: data_out = {8'd118, 8'd170, 1'b1, 1'b0};
5643: data_out = {8'd121, 8'd170, 1'b1, 1'b0};
5644: data_out = {8'd122, 8'd170, 1'b1, 1'b0};
5645: data_out = {8'd123, 8'd170, 1'b1, 1'b0};
5646: data_out = {8'd124, 8'd170, 1'b1, 1'b0};
5647: data_out = {8'd125, 8'd170, 1'b1, 1'b0};
5648: data_out = {8'd128, 8'd170, 1'b1, 1'b0};
5649: data_out = {8'd129, 8'd170, 1'b1, 1'b0};
5650: data_out = {8'd130, 8'd170, 1'b1, 1'b0};
5651: data_out = {8'd131, 8'd170, 1'b1, 1'b0};
5652: data_out = {8'd141, 8'd170, 1'b1, 1'b0};
5653: data_out = {8'd142, 8'd170, 1'b1, 1'b0};
5654: data_out = {8'd143, 8'd170, 1'b1, 1'b0};
5655: data_out = {8'd144, 8'd170, 1'b1, 1'b0};
5656: data_out = {8'd145, 8'd170, 1'b1, 1'b0};
5657: data_out = {8'd148, 8'd170, 1'b1, 1'b0};
5658: data_out = {8'd152, 8'd170, 1'b1, 1'b0};
5659: data_out = {8'd155, 8'd170, 1'b1, 1'b0};
5660: data_out = {8'd156, 8'd170, 1'b1, 1'b0};
5661: data_out = {8'd157, 8'd170, 1'b1, 1'b0};
5662: data_out = {8'd158, 8'd170, 1'b1, 1'b0};
5663: data_out = {8'd159, 8'd170, 1'b1, 1'b0};
5664: data_out = {8'd162, 8'd170, 1'b1, 1'b0};
5665: data_out = {8'd168, 8'd170, 1'b1, 1'b0};
5666: data_out = {8'd169, 8'd170, 1'b1, 1'b0};
5667: data_out = {8'd170, 8'd170, 1'b1, 1'b0};
5668: data_out = {8'd171, 8'd170, 1'b1, 1'b0};
5669: data_out = {8'd174, 8'd170, 1'b1, 1'b0};
5670: data_out = {8'd177, 8'd170, 1'b1, 1'b0};
5671: data_out = {8'd180, 8'd170, 1'b1, 1'b0};
5672: data_out = {8'd6, 8'd171, 1'b1, 1'b0};
5673: data_out = {8'd13, 8'd171, 1'b1, 1'b0};
5674: data_out = {8'd17, 8'd171, 1'b1, 1'b0};
5675: data_out = {8'd19, 8'd171, 1'b1, 1'b0};
5676: data_out = {8'd22, 8'd171, 1'b1, 1'b0};
5677: data_out = {8'd25, 8'd171, 1'b1, 1'b0};
5678: data_out = {8'd28, 8'd171, 1'b1, 1'b0};
5679: data_out = {8'd32, 8'd171, 1'b1, 1'b0};
5680: data_out = {8'd35, 8'd171, 1'b1, 1'b0};
5681: data_out = {8'd39, 8'd171, 1'b1, 1'b0};
5682: data_out = {8'd42, 8'd171, 1'b1, 1'b0};
5683: data_out = {8'd49, 8'd171, 1'b1, 1'b0};
5684: data_out = {8'd61, 8'd171, 1'b1, 1'b0};
5685: data_out = {8'd65, 8'd171, 1'b1, 1'b0};
5686: data_out = {8'd70, 8'd171, 1'b1, 1'b0};
5687: data_out = {8'd75, 8'd171, 1'b1, 1'b0};
5688: data_out = {8'd86, 8'd171, 1'b1, 1'b0};
5689: data_out = {8'd90, 8'd171, 1'b1, 1'b0};
5690: data_out = {8'd93, 8'd171, 1'b1, 1'b0};
5691: data_out = {8'd101, 8'd171, 1'b1, 1'b0};
5692: data_out = {8'd107, 8'd171, 1'b1, 1'b0};
5693: data_out = {8'd114, 8'd171, 1'b1, 1'b0};
5694: data_out = {8'd118, 8'd171, 1'b1, 1'b0};
5695: data_out = {8'd125, 8'd171, 1'b1, 1'b0};
5696: data_out = {8'd128, 8'd171, 1'b1, 1'b0};
5697: data_out = {8'd145, 8'd171, 1'b1, 1'b0};
5698: data_out = {8'd148, 8'd171, 1'b1, 1'b0};
5699: data_out = {8'd152, 8'd171, 1'b1, 1'b0};
5700: data_out = {8'd159, 8'd171, 1'b1, 1'b0};
5701: data_out = {8'd162, 8'd171, 1'b1, 1'b0};
5702: data_out = {8'd168, 8'd171, 1'b1, 1'b0};
5703: data_out = {8'd174, 8'd171, 1'b1, 1'b0};
5704: data_out = {8'd177, 8'd171, 1'b1, 1'b0};
5705: data_out = {8'd180, 8'd171, 1'b1, 1'b0};
5706: data_out = {8'd6, 8'd172, 1'b1, 1'b0};
5707: data_out = {8'd13, 8'd172, 1'b1, 1'b0};
5708: data_out = {8'd17, 8'd172, 1'b1, 1'b0};
5709: data_out = {8'd19, 8'd172, 1'b1, 1'b0};
5710: data_out = {8'd22, 8'd172, 1'b1, 1'b0};
5711: data_out = {8'd25, 8'd172, 1'b1, 1'b0};
5712: data_out = {8'd28, 8'd172, 1'b1, 1'b0};
5713: data_out = {8'd32, 8'd172, 1'b1, 1'b0};
5714: data_out = {8'd35, 8'd172, 1'b1, 1'b0};
5715: data_out = {8'd39, 8'd172, 1'b1, 1'b0};
5716: data_out = {8'd42, 8'd172, 1'b1, 1'b0};
5717: data_out = {8'd49, 8'd172, 1'b1, 1'b0};
5718: data_out = {8'd61, 8'd172, 1'b1, 1'b0};
5719: data_out = {8'd65, 8'd172, 1'b1, 1'b0};
5720: data_out = {8'd70, 8'd172, 1'b1, 1'b0};
5721: data_out = {8'd75, 8'd172, 1'b1, 1'b0};
5722: data_out = {8'd86, 8'd172, 1'b1, 1'b0};
5723: data_out = {8'd90, 8'd172, 1'b1, 1'b0};
5724: data_out = {8'd93, 8'd172, 1'b1, 1'b0};
5725: data_out = {8'd101, 8'd172, 1'b1, 1'b0};
5726: data_out = {8'd107, 8'd172, 1'b1, 1'b0};
5727: data_out = {8'd114, 8'd172, 1'b1, 1'b0};
5728: data_out = {8'd118, 8'd172, 1'b1, 1'b0};
5729: data_out = {8'd125, 8'd172, 1'b1, 1'b0};
5730: data_out = {8'd128, 8'd172, 1'b1, 1'b0};
5731: data_out = {8'd145, 8'd172, 1'b1, 1'b0};
5732: data_out = {8'd148, 8'd172, 1'b1, 1'b0};
5733: data_out = {8'd152, 8'd172, 1'b1, 1'b0};
5734: data_out = {8'd159, 8'd172, 1'b1, 1'b0};
5735: data_out = {8'd162, 8'd172, 1'b1, 1'b0};
5736: data_out = {8'd168, 8'd172, 1'b1, 1'b0};
5737: data_out = {8'd174, 8'd172, 1'b1, 1'b0};
5738: data_out = {8'd177, 8'd172, 1'b1, 1'b0};
5739: data_out = {8'd180, 8'd172, 1'b1, 1'b0};
5740: data_out = {8'd6, 8'd173, 1'b1, 1'b0};
5741: data_out = {8'd7, 8'd173, 1'b1, 1'b0};
5742: data_out = {8'd8, 8'd173, 1'b1, 1'b0};
5743: data_out = {8'd9, 8'd173, 1'b1, 1'b0};
5744: data_out = {8'd10, 8'd173, 1'b1, 1'b0};
5745: data_out = {8'd13, 8'd173, 1'b1, 1'b0};
5746: data_out = {8'd14, 8'd173, 1'b1, 1'b0};
5747: data_out = {8'd15, 8'd173, 1'b1, 1'b0};
5748: data_out = {8'd16, 8'd173, 1'b1, 1'b0};
5749: data_out = {8'd17, 8'd173, 1'b1, 1'b0};
5750: data_out = {8'd19, 8'd173, 1'b1, 1'b0};
5751: data_out = {8'd22, 8'd173, 1'b1, 1'b0};
5752: data_out = {8'd25, 8'd173, 1'b1, 1'b0};
5753: data_out = {8'd28, 8'd173, 1'b1, 1'b0};
5754: data_out = {8'd29, 8'd173, 1'b1, 1'b0};
5755: data_out = {8'd30, 8'd173, 1'b1, 1'b0};
5756: data_out = {8'd31, 8'd173, 1'b1, 1'b0};
5757: data_out = {8'd32, 8'd173, 1'b1, 1'b0};
5758: data_out = {8'd35, 8'd173, 1'b1, 1'b0};
5759: data_out = {8'd36, 8'd173, 1'b1, 1'b0};
5760: data_out = {8'd37, 8'd173, 1'b1, 1'b0};
5761: data_out = {8'd38, 8'd173, 1'b1, 1'b0};
5762: data_out = {8'd39, 8'd173, 1'b1, 1'b0};
5763: data_out = {8'd42, 8'd173, 1'b1, 1'b0};
5764: data_out = {8'd43, 8'd173, 1'b1, 1'b0};
5765: data_out = {8'd44, 8'd173, 1'b1, 1'b0};
5766: data_out = {8'd45, 8'd173, 1'b1, 1'b0};
5767: data_out = {8'd46, 8'd173, 1'b1, 1'b0};
5768: data_out = {8'd49, 8'd173, 1'b1, 1'b0};
5769: data_out = {8'd50, 8'd173, 1'b1, 1'b0};
5770: data_out = {8'd51, 8'd173, 1'b1, 1'b0};
5771: data_out = {8'd52, 8'd173, 1'b1, 1'b0};
5772: data_out = {8'd53, 8'd173, 1'b1, 1'b0};
5773: data_out = {8'd61, 8'd173, 1'b1, 1'b0};
5774: data_out = {8'd62, 8'd173, 1'b1, 1'b0};
5775: data_out = {8'd63, 8'd173, 1'b1, 1'b0};
5776: data_out = {8'd64, 8'd173, 1'b1, 1'b0};
5777: data_out = {8'd65, 8'd173, 1'b1, 1'b0};
5778: data_out = {8'd68, 8'd173, 1'b1, 1'b0};
5779: data_out = {8'd69, 8'd173, 1'b1, 1'b0};
5780: data_out = {8'd70, 8'd173, 1'b1, 1'b0};
5781: data_out = {8'd71, 8'd173, 1'b1, 1'b0};
5782: data_out = {8'd72, 8'd173, 1'b1, 1'b0};
5783: data_out = {8'd73, 8'd173, 1'b1, 1'b0};
5784: data_out = {8'd74, 8'd173, 1'b1, 1'b0};
5785: data_out = {8'd75, 8'd173, 1'b1, 1'b0};
5786: data_out = {8'd76, 8'd173, 1'b1, 1'b0};
5787: data_out = {8'd77, 8'd173, 1'b1, 1'b0};
5788: data_out = {8'd78, 8'd173, 1'b1, 1'b0};
5789: data_out = {8'd86, 8'd173, 1'b1, 1'b0};
5790: data_out = {8'd87, 8'd173, 1'b1, 1'b0};
5791: data_out = {8'd88, 8'd173, 1'b1, 1'b0};
5792: data_out = {8'd89, 8'd173, 1'b1, 1'b0};
5793: data_out = {8'd90, 8'd173, 1'b1, 1'b0};
5794: data_out = {8'd93, 8'd173, 1'b1, 1'b0};
5795: data_out = {8'd94, 8'd173, 1'b1, 1'b0};
5796: data_out = {8'd95, 8'd173, 1'b1, 1'b0};
5797: data_out = {8'd96, 8'd173, 1'b1, 1'b0};
5798: data_out = {8'd97, 8'd173, 1'b1, 1'b0};
5799: data_out = {8'd99, 8'd173, 1'b1, 1'b0};
5800: data_out = {8'd100, 8'd173, 1'b1, 1'b0};
5801: data_out = {8'd101, 8'd173, 1'b1, 1'b0};
5802: data_out = {8'd102, 8'd173, 1'b1, 1'b0};
5803: data_out = {8'd103, 8'd173, 1'b1, 1'b0};
5804: data_out = {8'd104, 8'd173, 1'b1, 1'b0};
5805: data_out = {8'd107, 8'd173, 1'b1, 1'b0};
5806: data_out = {8'd108, 8'd173, 1'b1, 1'b0};
5807: data_out = {8'd109, 8'd173, 1'b1, 1'b0};
5808: data_out = {8'd110, 8'd173, 1'b1, 1'b0};
5809: data_out = {8'd111, 8'd173, 1'b1, 1'b0};
5810: data_out = {8'd114, 8'd173, 1'b1, 1'b0};
5811: data_out = {8'd118, 8'd173, 1'b1, 1'b0};
5812: data_out = {8'd121, 8'd173, 1'b1, 1'b0};
5813: data_out = {8'd122, 8'd173, 1'b1, 1'b0};
5814: data_out = {8'd123, 8'd173, 1'b1, 1'b0};
5815: data_out = {8'd124, 8'd173, 1'b1, 1'b0};
5816: data_out = {8'd125, 8'd173, 1'b1, 1'b0};
5817: data_out = {8'd128, 8'd173, 1'b1, 1'b0};
5818: data_out = {8'd129, 8'd173, 1'b1, 1'b0};
5819: data_out = {8'd130, 8'd173, 1'b1, 1'b0};
5820: data_out = {8'd131, 8'd173, 1'b1, 1'b0};
5821: data_out = {8'd132, 8'd173, 1'b1, 1'b0};
5822: data_out = {8'd141, 8'd173, 1'b1, 1'b0};
5823: data_out = {8'd142, 8'd173, 1'b1, 1'b0};
5824: data_out = {8'd143, 8'd173, 1'b1, 1'b0};
5825: data_out = {8'd144, 8'd173, 1'b1, 1'b0};
5826: data_out = {8'd145, 8'd173, 1'b1, 1'b0};
5827: data_out = {8'd148, 8'd173, 1'b1, 1'b0};
5828: data_out = {8'd149, 8'd173, 1'b1, 1'b0};
5829: data_out = {8'd150, 8'd173, 1'b1, 1'b0};
5830: data_out = {8'd151, 8'd173, 1'b1, 1'b0};
5831: data_out = {8'd152, 8'd173, 1'b1, 1'b0};
5832: data_out = {8'd155, 8'd173, 1'b1, 1'b0};
5833: data_out = {8'd156, 8'd173, 1'b1, 1'b0};
5834: data_out = {8'd157, 8'd173, 1'b1, 1'b0};
5835: data_out = {8'd158, 8'd173, 1'b1, 1'b0};
5836: data_out = {8'd159, 8'd173, 1'b1, 1'b0};
5837: data_out = {8'd162, 8'd173, 1'b1, 1'b0};
5838: data_out = {8'd163, 8'd173, 1'b1, 1'b0};
5839: data_out = {8'd164, 8'd173, 1'b1, 1'b0};
5840: data_out = {8'd165, 8'd173, 1'b1, 1'b0};
5841: data_out = {8'd166, 8'd173, 1'b1, 1'b0};
5842: data_out = {8'd168, 8'd173, 1'b1, 1'b0};
5843: data_out = {8'd169, 8'd173, 1'b1, 1'b0};
5844: data_out = {8'd170, 8'd173, 1'b1, 1'b0};
5845: data_out = {8'd171, 8'd173, 1'b1, 1'b0};
5846: data_out = {8'd172, 8'd173, 1'b1, 1'b0};
5847: data_out = {8'd174, 8'd173, 1'b1, 1'b0};
5848: data_out = {8'd177, 8'd173, 1'b1, 1'b0};
5849: data_out = {8'd180, 8'd173, 1'b1, 1'b0};
5850: data_out = {8'd184, 8'd173, 1'b1, 1'b0};
5851: data_out = {8'd28, 8'd174, 1'b1, 1'b0};
5852: data_out = {8'd152, 8'd174, 1'b1, 1'b0};
5853: data_out = {8'd28, 8'd175, 1'b1, 1'b0};
5854: data_out = {8'd152, 8'd175, 1'b1, 1'b0};
5855: data_out = {8'd28, 8'd176, 1'b1, 1'b0};
5856: data_out = {8'd148, 8'd176, 1'b1, 1'b0};
5857: data_out = {8'd149, 8'd176, 1'b1, 1'b0};
5858: data_out = {8'd150, 8'd176, 1'b1, 1'b0};
5859: data_out = {8'd151, 8'd176, 1'b1, 1'b0};
5860: data_out = {8'd152, 8'd176, 1'b1, 1'b0};
5861: data_out = {8'd28, 8'd178, 1'b1, 1'b0};
5862: data_out = {8'd79, 8'd179, 1'b1, 1'b0};
5863: data_out = {8'd119, 8'd179, 1'b1, 1'b0};
5864: data_out = {8'd7, 8'd180, 1'b1, 1'b0};
5865: data_out = {8'd8, 8'd180, 1'b1, 1'b0};
5866: data_out = {8'd9, 8'd180, 1'b1, 1'b0};
5867: data_out = {8'd12, 8'd180, 1'b1, 1'b0};
5868: data_out = {8'd13, 8'd180, 1'b1, 1'b0};
5869: data_out = {8'd14, 8'd180, 1'b1, 1'b0};
5870: data_out = {8'd15, 8'd180, 1'b1, 1'b0};
5871: data_out = {8'd16, 8'd180, 1'b1, 1'b0};
5872: data_out = {8'd19, 8'd180, 1'b1, 1'b0};
5873: data_out = {8'd20, 8'd180, 1'b1, 1'b0};
5874: data_out = {8'd21, 8'd180, 1'b1, 1'b0};
5875: data_out = {8'd22, 8'd180, 1'b1, 1'b0};
5876: data_out = {8'd23, 8'd180, 1'b1, 1'b0};
5877: data_out = {8'd26, 8'd180, 1'b1, 1'b0};
5878: data_out = {8'd27, 8'd180, 1'b1, 1'b0};
5879: data_out = {8'd28, 8'd180, 1'b1, 1'b0};
5880: data_out = {8'd32, 8'd180, 1'b1, 1'b0};
5881: data_out = {8'd33, 8'd180, 1'b1, 1'b0};
5882: data_out = {8'd34, 8'd180, 1'b1, 1'b0};
5883: data_out = {8'd35, 8'd180, 1'b1, 1'b0};
5884: data_out = {8'd36, 8'd180, 1'b1, 1'b0};
5885: data_out = {8'd39, 8'd180, 1'b1, 1'b0};
5886: data_out = {8'd40, 8'd180, 1'b1, 1'b0};
5887: data_out = {8'd41, 8'd180, 1'b1, 1'b0};
5888: data_out = {8'd42, 8'd180, 1'b1, 1'b0};
5889: data_out = {8'd43, 8'd180, 1'b1, 1'b0};
5890: data_out = {8'd58, 8'd180, 1'b1, 1'b0};
5891: data_out = {8'd59, 8'd180, 1'b1, 1'b0};
5892: data_out = {8'd60, 8'd180, 1'b1, 1'b0};
5893: data_out = {8'd61, 8'd180, 1'b1, 1'b0};
5894: data_out = {8'd62, 8'd180, 1'b1, 1'b0};
5895: data_out = {8'd65, 8'd180, 1'b1, 1'b0};
5896: data_out = {8'd66, 8'd180, 1'b1, 1'b0};
5897: data_out = {8'd67, 8'd180, 1'b1, 1'b0};
5898: data_out = {8'd68, 8'd180, 1'b1, 1'b0};
5899: data_out = {8'd69, 8'd180, 1'b1, 1'b0};
5900: data_out = {8'd72, 8'd180, 1'b1, 1'b0};
5901: data_out = {8'd73, 8'd180, 1'b1, 1'b0};
5902: data_out = {8'd74, 8'd180, 1'b1, 1'b0};
5903: data_out = {8'd75, 8'd180, 1'b1, 1'b0};
5904: data_out = {8'd76, 8'd180, 1'b1, 1'b0};
5905: data_out = {8'd78, 8'd180, 1'b1, 1'b0};
5906: data_out = {8'd79, 8'd180, 1'b1, 1'b0};
5907: data_out = {8'd80, 8'd180, 1'b1, 1'b0};
5908: data_out = {8'd81, 8'd180, 1'b1, 1'b0};
5909: data_out = {8'd82, 8'd180, 1'b1, 1'b0};
5910: data_out = {8'd91, 8'd180, 1'b1, 1'b0};
5911: data_out = {8'd92, 8'd180, 1'b1, 1'b0};
5912: data_out = {8'd93, 8'd180, 1'b1, 1'b0};
5913: data_out = {8'd94, 8'd180, 1'b1, 1'b0};
5914: data_out = {8'd95, 8'd180, 1'b1, 1'b0};
5915: data_out = {8'd98, 8'd180, 1'b1, 1'b0};
5916: data_out = {8'd99, 8'd180, 1'b1, 1'b0};
5917: data_out = {8'd100, 8'd180, 1'b1, 1'b0};
5918: data_out = {8'd101, 8'd180, 1'b1, 1'b0};
5919: data_out = {8'd102, 8'd180, 1'b1, 1'b0};
5920: data_out = {8'd105, 8'd180, 1'b1, 1'b0};
5921: data_out = {8'd106, 8'd180, 1'b1, 1'b0};
5922: data_out = {8'd107, 8'd180, 1'b1, 1'b0};
5923: data_out = {8'd108, 8'd180, 1'b1, 1'b0};
5924: data_out = {8'd109, 8'd180, 1'b1, 1'b0};
5925: data_out = {8'd112, 8'd180, 1'b1, 1'b0};
5926: data_out = {8'd113, 8'd180, 1'b1, 1'b0};
5927: data_out = {8'd114, 8'd180, 1'b1, 1'b0};
5928: data_out = {8'd115, 8'd180, 1'b1, 1'b0};
5929: data_out = {8'd116, 8'd180, 1'b1, 1'b0};
5930: data_out = {8'd118, 8'd180, 1'b1, 1'b0};
5931: data_out = {8'd119, 8'd180, 1'b1, 1'b0};
5932: data_out = {8'd120, 8'd180, 1'b1, 1'b0};
5933: data_out = {8'd121, 8'd180, 1'b1, 1'b0};
5934: data_out = {8'd122, 8'd180, 1'b1, 1'b0};
5935: data_out = {8'd7, 8'd181, 1'b1, 1'b0};
5936: data_out = {8'd9, 8'd181, 1'b1, 1'b0};
5937: data_out = {8'd12, 8'd181, 1'b1, 1'b0};
5938: data_out = {8'd16, 8'd181, 1'b1, 1'b0};
5939: data_out = {8'd19, 8'd181, 1'b1, 1'b0};
5940: data_out = {8'd22, 8'd181, 1'b1, 1'b0};
5941: data_out = {8'd28, 8'd181, 1'b1, 1'b0};
5942: data_out = {8'd32, 8'd181, 1'b1, 1'b0};
5943: data_out = {8'd36, 8'd181, 1'b1, 1'b0};
5944: data_out = {8'd39, 8'd181, 1'b1, 1'b0};
5945: data_out = {8'd43, 8'd181, 1'b1, 1'b0};
5946: data_out = {8'd58, 8'd181, 1'b1, 1'b0};
5947: data_out = {8'd62, 8'd181, 1'b1, 1'b0};
5948: data_out = {8'd65, 8'd181, 1'b1, 1'b0};
5949: data_out = {8'd69, 8'd181, 1'b1, 1'b0};
5950: data_out = {8'd72, 8'd181, 1'b1, 1'b0};
5951: data_out = {8'd76, 8'd181, 1'b1, 1'b0};
5952: data_out = {8'd79, 8'd181, 1'b1, 1'b0};
5953: data_out = {8'd91, 8'd181, 1'b1, 1'b0};
5954: data_out = {8'd95, 8'd181, 1'b1, 1'b0};
5955: data_out = {8'd98, 8'd181, 1'b1, 1'b0};
5956: data_out = {8'd102, 8'd181, 1'b1, 1'b0};
5957: data_out = {8'd105, 8'd181, 1'b1, 1'b0};
5958: data_out = {8'd109, 8'd181, 1'b1, 1'b0};
5959: data_out = {8'd112, 8'd181, 1'b1, 1'b0};
5960: data_out = {8'd116, 8'd181, 1'b1, 1'b0};
5961: data_out = {8'd119, 8'd181, 1'b1, 1'b0};
5962: data_out = {8'd7, 8'd182, 1'b1, 1'b0};
5963: data_out = {8'd12, 8'd182, 1'b1, 1'b0};
5964: data_out = {8'd16, 8'd182, 1'b1, 1'b0};
5965: data_out = {8'd19, 8'd182, 1'b1, 1'b0};
5966: data_out = {8'd22, 8'd182, 1'b1, 1'b0};
5967: data_out = {8'd28, 8'd182, 1'b1, 1'b0};
5968: data_out = {8'd32, 8'd182, 1'b1, 1'b0};
5969: data_out = {8'd36, 8'd182, 1'b1, 1'b0};
5970: data_out = {8'd39, 8'd182, 1'b1, 1'b0};
5971: data_out = {8'd43, 8'd182, 1'b1, 1'b0};
5972: data_out = {8'd58, 8'd182, 1'b1, 1'b0};
5973: data_out = {8'd62, 8'd182, 1'b1, 1'b0};
5974: data_out = {8'd69, 8'd182, 1'b1, 1'b0};
5975: data_out = {8'd72, 8'd182, 1'b1, 1'b0};
5976: data_out = {8'd79, 8'd182, 1'b1, 1'b0};
5977: data_out = {8'd91, 8'd182, 1'b1, 1'b0};
5978: data_out = {8'd98, 8'd182, 1'b1, 1'b0};
5979: data_out = {8'd102, 8'd182, 1'b1, 1'b0};
5980: data_out = {8'd109, 8'd182, 1'b1, 1'b0};
5981: data_out = {8'd112, 8'd182, 1'b1, 1'b0};
5982: data_out = {8'd119, 8'd182, 1'b1, 1'b0};
5983: data_out = {8'd7, 8'd183, 1'b1, 1'b0};
5984: data_out = {8'd12, 8'd183, 1'b1, 1'b0};
5985: data_out = {8'd13, 8'd183, 1'b1, 1'b0};
5986: data_out = {8'd14, 8'd183, 1'b1, 1'b0};
5987: data_out = {8'd15, 8'd183, 1'b1, 1'b0};
5988: data_out = {8'd19, 8'd183, 1'b1, 1'b0};
5989: data_out = {8'd22, 8'd183, 1'b1, 1'b0};
5990: data_out = {8'd28, 8'd183, 1'b1, 1'b0};
5991: data_out = {8'd32, 8'd183, 1'b1, 1'b0};
5992: data_out = {8'd36, 8'd183, 1'b1, 1'b0};
5993: data_out = {8'd39, 8'd183, 1'b1, 1'b0};
5994: data_out = {8'd43, 8'd183, 1'b1, 1'b0};
5995: data_out = {8'd47, 8'd183, 1'b1, 1'b0};
5996: data_out = {8'd58, 8'd183, 1'b1, 1'b0};
5997: data_out = {8'd59, 8'd183, 1'b1, 1'b0};
5998: data_out = {8'd60, 8'd183, 1'b1, 1'b0};
5999: data_out = {8'd61, 8'd183, 1'b1, 1'b0};
6000: data_out = {8'd66, 8'd183, 1'b1, 1'b0};
6001: data_out = {8'd67, 8'd183, 1'b1, 1'b0};
6002: data_out = {8'd68, 8'd183, 1'b1, 1'b0};
6003: data_out = {8'd69, 8'd183, 1'b1, 1'b0};
6004: data_out = {8'd72, 8'd183, 1'b1, 1'b0};
6005: data_out = {8'd73, 8'd183, 1'b1, 1'b0};
6006: data_out = {8'd74, 8'd183, 1'b1, 1'b0};
6007: data_out = {8'd75, 8'd183, 1'b1, 1'b0};
6008: data_out = {8'd76, 8'd183, 1'b1, 1'b0};
6009: data_out = {8'd79, 8'd183, 1'b1, 1'b0};
6010: data_out = {8'd91, 8'd183, 1'b1, 1'b0};
6011: data_out = {8'd98, 8'd183, 1'b1, 1'b0};
6012: data_out = {8'd102, 8'd183, 1'b1, 1'b0};
6013: data_out = {8'd106, 8'd183, 1'b1, 1'b0};
6014: data_out = {8'd107, 8'd183, 1'b1, 1'b0};
6015: data_out = {8'd108, 8'd183, 1'b1, 1'b0};
6016: data_out = {8'd109, 8'd183, 1'b1, 1'b0};
6017: data_out = {8'd112, 8'd183, 1'b1, 1'b0};
6018: data_out = {8'd113, 8'd183, 1'b1, 1'b0};
6019: data_out = {8'd114, 8'd183, 1'b1, 1'b0};
6020: data_out = {8'd115, 8'd183, 1'b1, 1'b0};
6021: data_out = {8'd116, 8'd183, 1'b1, 1'b0};
6022: data_out = {8'd119, 8'd183, 1'b1, 1'b0};
6023: data_out = {8'd7, 8'd184, 1'b1, 1'b0};
6024: data_out = {8'd12, 8'd184, 1'b1, 1'b0};
6025: data_out = {8'd19, 8'd184, 1'b1, 1'b0};
6026: data_out = {8'd20, 8'd184, 1'b1, 1'b0};
6027: data_out = {8'd21, 8'd184, 1'b1, 1'b0};
6028: data_out = {8'd22, 8'd184, 1'b1, 1'b0};
6029: data_out = {8'd28, 8'd184, 1'b1, 1'b0};
6030: data_out = {8'd32, 8'd184, 1'b1, 1'b0};
6031: data_out = {8'd36, 8'd184, 1'b1, 1'b0};
6032: data_out = {8'd39, 8'd184, 1'b1, 1'b0};
6033: data_out = {8'd43, 8'd184, 1'b1, 1'b0};
6034: data_out = {8'd58, 8'd184, 1'b1, 1'b0};
6035: data_out = {8'd65, 8'd184, 1'b1, 1'b0};
6036: data_out = {8'd69, 8'd184, 1'b1, 1'b0};
6037: data_out = {8'd76, 8'd184, 1'b1, 1'b0};
6038: data_out = {8'd79, 8'd184, 1'b1, 1'b0};
6039: data_out = {8'd91, 8'd184, 1'b1, 1'b0};
6040: data_out = {8'd98, 8'd184, 1'b1, 1'b0};
6041: data_out = {8'd102, 8'd184, 1'b1, 1'b0};
6042: data_out = {8'd105, 8'd184, 1'b1, 1'b0};
6043: data_out = {8'd109, 8'd184, 1'b1, 1'b0};
6044: data_out = {8'd116, 8'd184, 1'b1, 1'b0};
6045: data_out = {8'd119, 8'd184, 1'b1, 1'b0};
6046: data_out = {8'd7, 8'd185, 1'b1, 1'b0};
6047: data_out = {8'd12, 8'd185, 1'b1, 1'b0};
6048: data_out = {8'd19, 8'd185, 1'b1, 1'b0};
6049: data_out = {8'd28, 8'd185, 1'b1, 1'b0};
6050: data_out = {8'd32, 8'd185, 1'b1, 1'b0};
6051: data_out = {8'd36, 8'd185, 1'b1, 1'b0};
6052: data_out = {8'd39, 8'd185, 1'b1, 1'b0};
6053: data_out = {8'd43, 8'd185, 1'b1, 1'b0};
6054: data_out = {8'd58, 8'd185, 1'b1, 1'b0};
6055: data_out = {8'd65, 8'd185, 1'b1, 1'b0};
6056: data_out = {8'd69, 8'd185, 1'b1, 1'b0};
6057: data_out = {8'd76, 8'd185, 1'b1, 1'b0};
6058: data_out = {8'd79, 8'd185, 1'b1, 1'b0};
6059: data_out = {8'd91, 8'd185, 1'b1, 1'b0};
6060: data_out = {8'd98, 8'd185, 1'b1, 1'b0};
6061: data_out = {8'd102, 8'd185, 1'b1, 1'b0};
6062: data_out = {8'd105, 8'd185, 1'b1, 1'b0};
6063: data_out = {8'd109, 8'd185, 1'b1, 1'b0};
6064: data_out = {8'd116, 8'd185, 1'b1, 1'b0};
6065: data_out = {8'd119, 8'd185, 1'b1, 1'b0};
6066: data_out = {8'd5, 8'd186, 1'b1, 1'b0};
6067: data_out = {8'd6, 8'd186, 1'b1, 1'b0};
6068: data_out = {8'd7, 8'd186, 1'b1, 1'b0};
6069: data_out = {8'd8, 8'd186, 1'b1, 1'b0};
6070: data_out = {8'd9, 8'd186, 1'b1, 1'b0};
6071: data_out = {8'd10, 8'd186, 1'b1, 1'b0};
6072: data_out = {8'd12, 8'd186, 1'b1, 1'b0};
6073: data_out = {8'd13, 8'd186, 1'b1, 1'b0};
6074: data_out = {8'd14, 8'd186, 1'b1, 1'b0};
6075: data_out = {8'd15, 8'd186, 1'b1, 1'b0};
6076: data_out = {8'd16, 8'd186, 1'b1, 1'b0};
6077: data_out = {8'd19, 8'd186, 1'b1, 1'b0};
6078: data_out = {8'd20, 8'd186, 1'b1, 1'b0};
6079: data_out = {8'd21, 8'd186, 1'b1, 1'b0};
6080: data_out = {8'd22, 8'd186, 1'b1, 1'b0};
6081: data_out = {8'd23, 8'd186, 1'b1, 1'b0};
6082: data_out = {8'd26, 8'd186, 1'b1, 1'b0};
6083: data_out = {8'd27, 8'd186, 1'b1, 1'b0};
6084: data_out = {8'd28, 8'd186, 1'b1, 1'b0};
6085: data_out = {8'd29, 8'd186, 1'b1, 1'b0};
6086: data_out = {8'd30, 8'd186, 1'b1, 1'b0};
6087: data_out = {8'd32, 8'd186, 1'b1, 1'b0};
6088: data_out = {8'd33, 8'd186, 1'b1, 1'b0};
6089: data_out = {8'd34, 8'd186, 1'b1, 1'b0};
6090: data_out = {8'd35, 8'd186, 1'b1, 1'b0};
6091: data_out = {8'd36, 8'd186, 1'b1, 1'b0};
6092: data_out = {8'd39, 8'd186, 1'b1, 1'b0};
6093: data_out = {8'd43, 8'd186, 1'b1, 1'b0};
6094: data_out = {8'd47, 8'd186, 1'b1, 1'b0};
6095: data_out = {8'd58, 8'd186, 1'b1, 1'b0};
6096: data_out = {8'd59, 8'd186, 1'b1, 1'b0};
6097: data_out = {8'd60, 8'd186, 1'b1, 1'b0};
6098: data_out = {8'd61, 8'd186, 1'b1, 1'b0};
6099: data_out = {8'd62, 8'd186, 1'b1, 1'b0};
6100: data_out = {8'd65, 8'd186, 1'b1, 1'b0};
6101: data_out = {8'd66, 8'd186, 1'b1, 1'b0};
6102: data_out = {8'd67, 8'd186, 1'b1, 1'b0};
6103: data_out = {8'd68, 8'd186, 1'b1, 1'b0};
6104: data_out = {8'd69, 8'd186, 1'b1, 1'b0};
6105: data_out = {8'd72, 8'd186, 1'b1, 1'b0};
6106: data_out = {8'd73, 8'd186, 1'b1, 1'b0};
6107: data_out = {8'd74, 8'd186, 1'b1, 1'b0};
6108: data_out = {8'd75, 8'd186, 1'b1, 1'b0};
6109: data_out = {8'd76, 8'd186, 1'b1, 1'b0};
6110: data_out = {8'd79, 8'd186, 1'b1, 1'b0};
6111: data_out = {8'd80, 8'd186, 1'b1, 1'b0};
6112: data_out = {8'd81, 8'd186, 1'b1, 1'b0};
6113: data_out = {8'd82, 8'd186, 1'b1, 1'b0};
6114: data_out = {8'd83, 8'd186, 1'b1, 1'b0};
6115: data_out = {8'd91, 8'd186, 1'b1, 1'b0};
6116: data_out = {8'd92, 8'd186, 1'b1, 1'b0};
6117: data_out = {8'd93, 8'd186, 1'b1, 1'b0};
6118: data_out = {8'd94, 8'd186, 1'b1, 1'b0};
6119: data_out = {8'd95, 8'd186, 1'b1, 1'b0};
6120: data_out = {8'd98, 8'd186, 1'b1, 1'b0};
6121: data_out = {8'd99, 8'd186, 1'b1, 1'b0};
6122: data_out = {8'd100, 8'd186, 1'b1, 1'b0};
6123: data_out = {8'd101, 8'd186, 1'b1, 1'b0};
6124: data_out = {8'd102, 8'd186, 1'b1, 1'b0};
6125: data_out = {8'd105, 8'd186, 1'b1, 1'b0};
6126: data_out = {8'd106, 8'd186, 1'b1, 1'b0};
6127: data_out = {8'd107, 8'd186, 1'b1, 1'b0};
6128: data_out = {8'd108, 8'd186, 1'b1, 1'b0};
6129: data_out = {8'd109, 8'd186, 1'b1, 1'b0};
6130: data_out = {8'd112, 8'd186, 1'b1, 1'b0};
6131: data_out = {8'd113, 8'd186, 1'b1, 1'b0};
6132: data_out = {8'd114, 8'd186, 1'b1, 1'b0};
6133: data_out = {8'd115, 8'd186, 1'b1, 1'b0};
6134: data_out = {8'd116, 8'd186, 1'b1, 1'b0};
6135: data_out = {8'd119, 8'd186, 1'b1, 1'b0};
6136: data_out = {8'd120, 8'd186, 1'b1, 1'b0};
6137: data_out = {8'd121, 8'd186, 1'b1, 1'b0};
6138: data_out = {8'd122, 8'd186, 1'b1, 1'b0};
6139: data_out = {8'd123, 8'd186, 1'b1, 1'b0};
6140: data_out = {8'd19, 8'd187, 1'b1, 1'b0};
6141: data_out = {8'd23, 8'd187, 1'b1, 1'b0};
6142: data_out = {8'd19, 8'd188, 1'b1, 1'b0};
6143: data_out = {8'd23, 8'd188, 1'b1, 1'b0};
6144: data_out = {8'd19, 8'd189, 1'b1, 1'b0};
6145: data_out = {8'd20, 8'd189, 1'b1, 1'b0};
6146: data_out = {8'd21, 8'd189, 1'b1, 1'b0};
6147: data_out = {8'd22, 8'd189, 1'b1, 1'b0};
6148: data_out = {8'd23, 8'd189, 1'b1, 1'b0};
6149: data_out = {8'd89, 8'd191, 1'b1, 1'b0};
6150: data_out = {8'd92, 8'd191, 1'b1, 1'b0};
6151: data_out = {8'd13, 8'd192, 1'b1, 1'b0};
6152: data_out = {8'd26, 8'd192, 1'b1, 1'b0};
6153: data_out = {8'd65, 8'd192, 1'b1, 1'b0};
6154: data_out = {8'd89, 8'd192, 1'b1, 1'b0};
6155: data_out = {8'd92, 8'd192, 1'b1, 1'b0};
6156: data_out = {8'd6, 8'd193, 1'b1, 1'b0};
6157: data_out = {8'd7, 8'd193, 1'b1, 1'b0};
6158: data_out = {8'd8, 8'd193, 1'b1, 1'b0};
6159: data_out = {8'd9, 8'd193, 1'b1, 1'b0};
6160: data_out = {8'd10, 8'd193, 1'b1, 1'b0};
6161: data_out = {8'd12, 8'd193, 1'b1, 1'b0};
6162: data_out = {8'd13, 8'd193, 1'b1, 1'b0};
6163: data_out = {8'd14, 8'd193, 1'b1, 1'b0};
6164: data_out = {8'd15, 8'd193, 1'b1, 1'b0};
6165: data_out = {8'd16, 8'd193, 1'b1, 1'b0};
6166: data_out = {8'd19, 8'd193, 1'b1, 1'b0};
6167: data_out = {8'd20, 8'd193, 1'b1, 1'b0};
6168: data_out = {8'd21, 8'd193, 1'b1, 1'b0};
6169: data_out = {8'd22, 8'd193, 1'b1, 1'b0};
6170: data_out = {8'd23, 8'd193, 1'b1, 1'b0};
6171: data_out = {8'd25, 8'd193, 1'b1, 1'b0};
6172: data_out = {8'd26, 8'd193, 1'b1, 1'b0};
6173: data_out = {8'd27, 8'd193, 1'b1, 1'b0};
6174: data_out = {8'd28, 8'd193, 1'b1, 1'b0};
6175: data_out = {8'd29, 8'd193, 1'b1, 1'b0};
6176: data_out = {8'd32, 8'd193, 1'b1, 1'b0};
6177: data_out = {8'd36, 8'd193, 1'b1, 1'b0};
6178: data_out = {8'd39, 8'd193, 1'b1, 1'b0};
6179: data_out = {8'd40, 8'd193, 1'b1, 1'b0};
6180: data_out = {8'd41, 8'd193, 1'b1, 1'b0};
6181: data_out = {8'd42, 8'd193, 1'b1, 1'b0};
6182: data_out = {8'd43, 8'd193, 1'b1, 1'b0};
6183: data_out = {8'd58, 8'd193, 1'b1, 1'b0};
6184: data_out = {8'd59, 8'd193, 1'b1, 1'b0};
6185: data_out = {8'd60, 8'd193, 1'b1, 1'b0};
6186: data_out = {8'd61, 8'd193, 1'b1, 1'b0};
6187: data_out = {8'd62, 8'd193, 1'b1, 1'b0};
6188: data_out = {8'd64, 8'd193, 1'b1, 1'b0};
6189: data_out = {8'd65, 8'd193, 1'b1, 1'b0};
6190: data_out = {8'd66, 8'd193, 1'b1, 1'b0};
6191: data_out = {8'd67, 8'd193, 1'b1, 1'b0};
6192: data_out = {8'd68, 8'd193, 1'b1, 1'b0};
6193: data_out = {8'd71, 8'd193, 1'b1, 1'b0};
6194: data_out = {8'd72, 8'd193, 1'b1, 1'b0};
6195: data_out = {8'd73, 8'd193, 1'b1, 1'b0};
6196: data_out = {8'd74, 8'd193, 1'b1, 1'b0};
6197: data_out = {8'd75, 8'd193, 1'b1, 1'b0};
6198: data_out = {8'd78, 8'd193, 1'b1, 1'b0};
6199: data_out = {8'd79, 8'd193, 1'b1, 1'b0};
6200: data_out = {8'd80, 8'd193, 1'b1, 1'b0};
6201: data_out = {8'd81, 8'd193, 1'b1, 1'b0};
6202: data_out = {8'd82, 8'd193, 1'b1, 1'b0};
6203: data_out = {8'd85, 8'd193, 1'b1, 1'b0};
6204: data_out = {8'd86, 8'd193, 1'b1, 1'b0};
6205: data_out = {8'd87, 8'd193, 1'b1, 1'b0};
6206: data_out = {8'd88, 8'd193, 1'b1, 1'b0};
6207: data_out = {8'd89, 8'd193, 1'b1, 1'b0};
6208: data_out = {8'd92, 8'd193, 1'b1, 1'b0};
6209: data_out = {8'd93, 8'd193, 1'b1, 1'b0};
6210: data_out = {8'd94, 8'd193, 1'b1, 1'b0};
6211: data_out = {8'd95, 8'd193, 1'b1, 1'b0};
6212: data_out = {8'd96, 8'd193, 1'b1, 1'b0};
6213: data_out = {8'd99, 8'd193, 1'b1, 1'b0};
6214: data_out = {8'd103, 8'd193, 1'b1, 1'b0};
6215: data_out = {8'd6, 8'd194, 1'b1, 1'b0};
6216: data_out = {8'd10, 8'd194, 1'b1, 1'b0};
6217: data_out = {8'd13, 8'd194, 1'b1, 1'b0};
6218: data_out = {8'd19, 8'd194, 1'b1, 1'b0};
6219: data_out = {8'd23, 8'd194, 1'b1, 1'b0};
6220: data_out = {8'd26, 8'd194, 1'b1, 1'b0};
6221: data_out = {8'd32, 8'd194, 1'b1, 1'b0};
6222: data_out = {8'd36, 8'd194, 1'b1, 1'b0};
6223: data_out = {8'd39, 8'd194, 1'b1, 1'b0};
6224: data_out = {8'd43, 8'd194, 1'b1, 1'b0};
6225: data_out = {8'd58, 8'd194, 1'b1, 1'b0};
6226: data_out = {8'd62, 8'd194, 1'b1, 1'b0};
6227: data_out = {8'd65, 8'd194, 1'b1, 1'b0};
6228: data_out = {8'd71, 8'd194, 1'b1, 1'b0};
6229: data_out = {8'd75, 8'd194, 1'b1, 1'b0};
6230: data_out = {8'd78, 8'd194, 1'b1, 1'b0};
6231: data_out = {8'd82, 8'd194, 1'b1, 1'b0};
6232: data_out = {8'd85, 8'd194, 1'b1, 1'b0};
6233: data_out = {8'd89, 8'd194, 1'b1, 1'b0};
6234: data_out = {8'd92, 8'd194, 1'b1, 1'b0};
6235: data_out = {8'd96, 8'd194, 1'b1, 1'b0};
6236: data_out = {8'd99, 8'd194, 1'b1, 1'b0};
6237: data_out = {8'd103, 8'd194, 1'b1, 1'b0};
6238: data_out = {8'd6, 8'd195, 1'b1, 1'b0};
6239: data_out = {8'd13, 8'd195, 1'b1, 1'b0};
6240: data_out = {8'd23, 8'd195, 1'b1, 1'b0};
6241: data_out = {8'd26, 8'd195, 1'b1, 1'b0};
6242: data_out = {8'd32, 8'd195, 1'b1, 1'b0};
6243: data_out = {8'd36, 8'd195, 1'b1, 1'b0};
6244: data_out = {8'd39, 8'd195, 1'b1, 1'b0};
6245: data_out = {8'd58, 8'd195, 1'b1, 1'b0};
6246: data_out = {8'd65, 8'd195, 1'b1, 1'b0};
6247: data_out = {8'd75, 8'd195, 1'b1, 1'b0};
6248: data_out = {8'd78, 8'd195, 1'b1, 1'b0};
6249: data_out = {8'd82, 8'd195, 1'b1, 1'b0};
6250: data_out = {8'd85, 8'd195, 1'b1, 1'b0};
6251: data_out = {8'd89, 8'd195, 1'b1, 1'b0};
6252: data_out = {8'd92, 8'd195, 1'b1, 1'b0};
6253: data_out = {8'd96, 8'd195, 1'b1, 1'b0};
6254: data_out = {8'd99, 8'd195, 1'b1, 1'b0};
6255: data_out = {8'd103, 8'd195, 1'b1, 1'b0};
6256: data_out = {8'd6, 8'd196, 1'b1, 1'b0};
6257: data_out = {8'd7, 8'd196, 1'b1, 1'b0};
6258: data_out = {8'd8, 8'd196, 1'b1, 1'b0};
6259: data_out = {8'd9, 8'd196, 1'b1, 1'b0};
6260: data_out = {8'd10, 8'd196, 1'b1, 1'b0};
6261: data_out = {8'd13, 8'd196, 1'b1, 1'b0};
6262: data_out = {8'd20, 8'd196, 1'b1, 1'b0};
6263: data_out = {8'd21, 8'd196, 1'b1, 1'b0};
6264: data_out = {8'd22, 8'd196, 1'b1, 1'b0};
6265: data_out = {8'd23, 8'd196, 1'b1, 1'b0};
6266: data_out = {8'd26, 8'd196, 1'b1, 1'b0};
6267: data_out = {8'd32, 8'd196, 1'b1, 1'b0};
6268: data_out = {8'd36, 8'd196, 1'b1, 1'b0};
6269: data_out = {8'd39, 8'd196, 1'b1, 1'b0};
6270: data_out = {8'd40, 8'd196, 1'b1, 1'b0};
6271: data_out = {8'd41, 8'd196, 1'b1, 1'b0};
6272: data_out = {8'd42, 8'd196, 1'b1, 1'b0};
6273: data_out = {8'd43, 8'd196, 1'b1, 1'b0};
6274: data_out = {8'd47, 8'd196, 1'b1, 1'b0};
6275: data_out = {8'd58, 8'd196, 1'b1, 1'b0};
6276: data_out = {8'd59, 8'd196, 1'b1, 1'b0};
6277: data_out = {8'd60, 8'd196, 1'b1, 1'b0};
6278: data_out = {8'd61, 8'd196, 1'b1, 1'b0};
6279: data_out = {8'd62, 8'd196, 1'b1, 1'b0};
6280: data_out = {8'd65, 8'd196, 1'b1, 1'b0};
6281: data_out = {8'd72, 8'd196, 1'b1, 1'b0};
6282: data_out = {8'd73, 8'd196, 1'b1, 1'b0};
6283: data_out = {8'd74, 8'd196, 1'b1, 1'b0};
6284: data_out = {8'd75, 8'd196, 1'b1, 1'b0};
6285: data_out = {8'd78, 8'd196, 1'b1, 1'b0};
6286: data_out = {8'd82, 8'd196, 1'b1, 1'b0};
6287: data_out = {8'd85, 8'd196, 1'b1, 1'b0};
6288: data_out = {8'd89, 8'd196, 1'b1, 1'b0};
6289: data_out = {8'd92, 8'd196, 1'b1, 1'b0};
6290: data_out = {8'd96, 8'd196, 1'b1, 1'b0};
6291: data_out = {8'd99, 8'd196, 1'b1, 1'b0};
6292: data_out = {8'd103, 8'd196, 1'b1, 1'b0};
6293: data_out = {8'd10, 8'd197, 1'b1, 1'b0};
6294: data_out = {8'd13, 8'd197, 1'b1, 1'b0};
6295: data_out = {8'd19, 8'd197, 1'b1, 1'b0};
6296: data_out = {8'd23, 8'd197, 1'b1, 1'b0};
6297: data_out = {8'd26, 8'd197, 1'b1, 1'b0};
6298: data_out = {8'd32, 8'd197, 1'b1, 1'b0};
6299: data_out = {8'd36, 8'd197, 1'b1, 1'b0};
6300: data_out = {8'd43, 8'd197, 1'b1, 1'b0};
6301: data_out = {8'd62, 8'd197, 1'b1, 1'b0};
6302: data_out = {8'd65, 8'd197, 1'b1, 1'b0};
6303: data_out = {8'd71, 8'd197, 1'b1, 1'b0};
6304: data_out = {8'd75, 8'd197, 1'b1, 1'b0};
6305: data_out = {8'd78, 8'd197, 1'b1, 1'b0};
6306: data_out = {8'd82, 8'd197, 1'b1, 1'b0};
6307: data_out = {8'd85, 8'd197, 1'b1, 1'b0};
6308: data_out = {8'd89, 8'd197, 1'b1, 1'b0};
6309: data_out = {8'd92, 8'd197, 1'b1, 1'b0};
6310: data_out = {8'd96, 8'd197, 1'b1, 1'b0};
6311: data_out = {8'd99, 8'd197, 1'b1, 1'b0};
6312: data_out = {8'd103, 8'd197, 1'b1, 1'b0};
6313: data_out = {8'd10, 8'd198, 1'b1, 1'b0};
6314: data_out = {8'd13, 8'd198, 1'b1, 1'b0};
6315: data_out = {8'd19, 8'd198, 1'b1, 1'b0};
6316: data_out = {8'd23, 8'd198, 1'b1, 1'b0};
6317: data_out = {8'd26, 8'd198, 1'b1, 1'b0};
6318: data_out = {8'd32, 8'd198, 1'b1, 1'b0};
6319: data_out = {8'd36, 8'd198, 1'b1, 1'b0};
6320: data_out = {8'd43, 8'd198, 1'b1, 1'b0};
6321: data_out = {8'd62, 8'd198, 1'b1, 1'b0};
6322: data_out = {8'd65, 8'd198, 1'b1, 1'b0};
6323: data_out = {8'd71, 8'd198, 1'b1, 1'b0};
6324: data_out = {8'd75, 8'd198, 1'b1, 1'b0};
6325: data_out = {8'd78, 8'd198, 1'b1, 1'b0};
6326: data_out = {8'd82, 8'd198, 1'b1, 1'b0};
6327: data_out = {8'd85, 8'd198, 1'b1, 1'b0};
6328: data_out = {8'd89, 8'd198, 1'b1, 1'b0};
6329: data_out = {8'd92, 8'd198, 1'b1, 1'b0};
6330: data_out = {8'd96, 8'd198, 1'b1, 1'b0};
6331: data_out = {8'd99, 8'd198, 1'b1, 1'b0};
6332: data_out = {8'd103, 8'd198, 1'b1, 1'b0};
6333: data_out = {8'd6, 8'd199, 1'b1, 1'b0};
6334: data_out = {8'd7, 8'd199, 1'b1, 1'b0};
6335: data_out = {8'd8, 8'd199, 1'b1, 1'b0};
6336: data_out = {8'd9, 8'd199, 1'b1, 1'b0};
6337: data_out = {8'd10, 8'd199, 1'b1, 1'b0};
6338: data_out = {8'd13, 8'd199, 1'b1, 1'b0};
6339: data_out = {8'd14, 8'd199, 1'b1, 1'b0};
6340: data_out = {8'd15, 8'd199, 1'b1, 1'b0};
6341: data_out = {8'd16, 8'd199, 1'b1, 1'b0};
6342: data_out = {8'd17, 8'd199, 1'b1, 1'b0};
6343: data_out = {8'd19, 8'd199, 1'b1, 1'b0};
6344: data_out = {8'd20, 8'd199, 1'b1, 1'b0};
6345: data_out = {8'd21, 8'd199, 1'b1, 1'b0};
6346: data_out = {8'd22, 8'd199, 1'b1, 1'b0};
6347: data_out = {8'd23, 8'd199, 1'b1, 1'b0};
6348: data_out = {8'd26, 8'd199, 1'b1, 1'b0};
6349: data_out = {8'd27, 8'd199, 1'b1, 1'b0};
6350: data_out = {8'd28, 8'd199, 1'b1, 1'b0};
6351: data_out = {8'd29, 8'd199, 1'b1, 1'b0};
6352: data_out = {8'd30, 8'd199, 1'b1, 1'b0};
6353: data_out = {8'd32, 8'd199, 1'b1, 1'b0};
6354: data_out = {8'd33, 8'd199, 1'b1, 1'b0};
6355: data_out = {8'd34, 8'd199, 1'b1, 1'b0};
6356: data_out = {8'd35, 8'd199, 1'b1, 1'b0};
6357: data_out = {8'd36, 8'd199, 1'b1, 1'b0};
6358: data_out = {8'd39, 8'd199, 1'b1, 1'b0};
6359: data_out = {8'd40, 8'd199, 1'b1, 1'b0};
6360: data_out = {8'd41, 8'd199, 1'b1, 1'b0};
6361: data_out = {8'd42, 8'd199, 1'b1, 1'b0};
6362: data_out = {8'd43, 8'd199, 1'b1, 1'b0};
6363: data_out = {8'd47, 8'd199, 1'b1, 1'b0};
6364: data_out = {8'd58, 8'd199, 1'b1, 1'b0};
6365: data_out = {8'd59, 8'd199, 1'b1, 1'b0};
6366: data_out = {8'd60, 8'd199, 1'b1, 1'b0};
6367: data_out = {8'd61, 8'd199, 1'b1, 1'b0};
6368: data_out = {8'd62, 8'd199, 1'b1, 1'b0};
6369: data_out = {8'd65, 8'd199, 1'b1, 1'b0};
6370: data_out = {8'd66, 8'd199, 1'b1, 1'b0};
6371: data_out = {8'd67, 8'd199, 1'b1, 1'b0};
6372: data_out = {8'd68, 8'd199, 1'b1, 1'b0};
6373: data_out = {8'd69, 8'd199, 1'b1, 1'b0};
6374: data_out = {8'd71, 8'd199, 1'b1, 1'b0};
6375: data_out = {8'd72, 8'd199, 1'b1, 1'b0};
6376: data_out = {8'd73, 8'd199, 1'b1, 1'b0};
6377: data_out = {8'd74, 8'd199, 1'b1, 1'b0};
6378: data_out = {8'd75, 8'd199, 1'b1, 1'b0};
6379: data_out = {8'd78, 8'd199, 1'b1, 1'b0};
6380: data_out = {8'd82, 8'd199, 1'b1, 1'b0};
6381: data_out = {8'd85, 8'd199, 1'b1, 1'b0};
6382: data_out = {8'd86, 8'd199, 1'b1, 1'b0};
6383: data_out = {8'd87, 8'd199, 1'b1, 1'b0};
6384: data_out = {8'd88, 8'd199, 1'b1, 1'b0};
6385: data_out = {8'd89, 8'd199, 1'b1, 1'b0};
6386: data_out = {8'd92, 8'd199, 1'b1, 1'b0};
6387: data_out = {8'd93, 8'd199, 1'b1, 1'b0};
6388: data_out = {8'd94, 8'd199, 1'b1, 1'b0};
6389: data_out = {8'd95, 8'd199, 1'b1, 1'b0};
6390: data_out = {8'd96, 8'd199, 1'b1, 1'b0};
6391: data_out = {8'd99, 8'd199, 1'b1, 1'b0};
6392: data_out = {8'd100, 8'd199, 1'b1, 1'b0};
6393: data_out = {8'd101, 8'd199, 1'b1, 1'b0};
6394: data_out = {8'd102, 8'd199, 1'b1, 1'b0};
6395: data_out = {8'd103, 8'd199, 1'b1, 1'b0};
6396: data_out = {8'd103, 8'd200, 1'b1, 1'b0};
6397: data_out = {8'd103, 8'd201, 1'b1, 1'b0};
6398: data_out = {8'd99, 8'd202, 1'b1, 1'b0};
6399: data_out = {8'd100, 8'd202, 1'b1, 1'b0};
6400: data_out = {8'd101, 8'd202, 1'b1, 1'b0};
6401: data_out = {8'd102, 8'd202, 1'b1, 1'b0};
6402: data_out = {8'd103, 8'd202, 1'b1, 1'b0};
6403: data_out = {8'd25, 8'd204, 1'b1, 1'b0};
6404: data_out = {8'd35, 8'd204, 1'b1, 1'b0};
6405: data_out = {8'd36, 8'd204, 1'b1, 1'b0};
6406: data_out = {8'd37, 8'd204, 1'b1, 1'b0};
6407: data_out = {8'd75, 8'd204, 1'b1, 1'b0};
6408: data_out = {8'd76, 8'd204, 1'b1, 1'b0};
6409: data_out = {8'd77, 8'd204, 1'b1, 1'b0};
6410: data_out = {8'd83, 8'd204, 1'b1, 1'b0};
6411: data_out = {8'd130, 8'd204, 1'b1, 1'b0};
6412: data_out = {8'd25, 8'd205, 1'b1, 1'b0};
6413: data_out = {8'd37, 8'd205, 1'b1, 1'b0};
6414: data_out = {8'd77, 8'd205, 1'b1, 1'b0};
6415: data_out = {8'd130, 8'd205, 1'b1, 1'b0};
6416: data_out = {8'd5, 8'd206, 1'b1, 1'b0};
6417: data_out = {8'd6, 8'd206, 1'b1, 1'b0};
6418: data_out = {8'd7, 8'd206, 1'b1, 1'b0};
6419: data_out = {8'd8, 8'd206, 1'b1, 1'b0};
6420: data_out = {8'd9, 8'd206, 1'b1, 1'b0};
6421: data_out = {8'd10, 8'd206, 1'b1, 1'b0};
6422: data_out = {8'd11, 8'd206, 1'b1, 1'b0};
6423: data_out = {8'd14, 8'd206, 1'b1, 1'b0};
6424: data_out = {8'd15, 8'd206, 1'b1, 1'b0};
6425: data_out = {8'd16, 8'd206, 1'b1, 1'b0};
6426: data_out = {8'd17, 8'd206, 1'b1, 1'b0};
6427: data_out = {8'd18, 8'd206, 1'b1, 1'b0};
6428: data_out = {8'd21, 8'd206, 1'b1, 1'b0};
6429: data_out = {8'd22, 8'd206, 1'b1, 1'b0};
6430: data_out = {8'd23, 8'd206, 1'b1, 1'b0};
6431: data_out = {8'd24, 8'd206, 1'b1, 1'b0};
6432: data_out = {8'd25, 8'd206, 1'b1, 1'b0};
6433: data_out = {8'd28, 8'd206, 1'b1, 1'b0};
6434: data_out = {8'd32, 8'd206, 1'b1, 1'b0};
6435: data_out = {8'd37, 8'd206, 1'b1, 1'b0};
6436: data_out = {8'd41, 8'd206, 1'b1, 1'b0};
6437: data_out = {8'd42, 8'd206, 1'b1, 1'b0};
6438: data_out = {8'd43, 8'd206, 1'b1, 1'b0};
6439: data_out = {8'd44, 8'd206, 1'b1, 1'b0};
6440: data_out = {8'd45, 8'd206, 1'b1, 1'b0};
6441: data_out = {8'd48, 8'd206, 1'b1, 1'b0};
6442: data_out = {8'd49, 8'd206, 1'b1, 1'b0};
6443: data_out = {8'd50, 8'd206, 1'b1, 1'b0};
6444: data_out = {8'd51, 8'd206, 1'b1, 1'b0};
6445: data_out = {8'd52, 8'd206, 1'b1, 1'b0};
6446: data_out = {8'd61, 8'd206, 1'b1, 1'b0};
6447: data_out = {8'd62, 8'd206, 1'b1, 1'b0};
6448: data_out = {8'd63, 8'd206, 1'b1, 1'b0};
6449: data_out = {8'd64, 8'd206, 1'b1, 1'b0};
6450: data_out = {8'd65, 8'd206, 1'b1, 1'b0};
6451: data_out = {8'd68, 8'd206, 1'b1, 1'b0};
6452: data_out = {8'd69, 8'd206, 1'b1, 1'b0};
6453: data_out = {8'd70, 8'd206, 1'b1, 1'b0};
6454: data_out = {8'd71, 8'd206, 1'b1, 1'b0};
6455: data_out = {8'd72, 8'd206, 1'b1, 1'b0};
6456: data_out = {8'd77, 8'd206, 1'b1, 1'b0};
6457: data_out = {8'd81, 8'd206, 1'b1, 1'b0};
6458: data_out = {8'd82, 8'd206, 1'b1, 1'b0};
6459: data_out = {8'd83, 8'd206, 1'b1, 1'b0};
6460: data_out = {8'd87, 8'd206, 1'b1, 1'b0};
6461: data_out = {8'd88, 8'd206, 1'b1, 1'b0};
6462: data_out = {8'd89, 8'd206, 1'b1, 1'b0};
6463: data_out = {8'd90, 8'd206, 1'b1, 1'b0};
6464: data_out = {8'd91, 8'd206, 1'b1, 1'b0};
6465: data_out = {8'd94, 8'd206, 1'b1, 1'b0};
6466: data_out = {8'd95, 8'd206, 1'b1, 1'b0};
6467: data_out = {8'd96, 8'd206, 1'b1, 1'b0};
6468: data_out = {8'd97, 8'd206, 1'b1, 1'b0};
6469: data_out = {8'd98, 8'd206, 1'b1, 1'b0};
6470: data_out = {8'd114, 8'd206, 1'b1, 1'b0};
6471: data_out = {8'd115, 8'd206, 1'b1, 1'b0};
6472: data_out = {8'd116, 8'd206, 1'b1, 1'b0};
6473: data_out = {8'd119, 8'd206, 1'b1, 1'b0};
6474: data_out = {8'd120, 8'd206, 1'b1, 1'b0};
6475: data_out = {8'd121, 8'd206, 1'b1, 1'b0};
6476: data_out = {8'd122, 8'd206, 1'b1, 1'b0};
6477: data_out = {8'd123, 8'd206, 1'b1, 1'b0};
6478: data_out = {8'd126, 8'd206, 1'b1, 1'b0};
6479: data_out = {8'd127, 8'd206, 1'b1, 1'b0};
6480: data_out = {8'd128, 8'd206, 1'b1, 1'b0};
6481: data_out = {8'd129, 8'd206, 1'b1, 1'b0};
6482: data_out = {8'd130, 8'd206, 1'b1, 1'b0};
6483: data_out = {8'd133, 8'd206, 1'b1, 1'b0};
6484: data_out = {8'd134, 8'd206, 1'b1, 1'b0};
6485: data_out = {8'd135, 8'd206, 1'b1, 1'b0};
6486: data_out = {8'd136, 8'd206, 1'b1, 1'b0};
6487: data_out = {8'd137, 8'd206, 1'b1, 1'b0};
6488: data_out = {8'd141, 8'd206, 1'b1, 1'b0};
6489: data_out = {8'd142, 8'd206, 1'b1, 1'b0};
6490: data_out = {8'd143, 8'd206, 1'b1, 1'b0};
6491: data_out = {8'd5, 8'd207, 1'b1, 1'b0};
6492: data_out = {8'd8, 8'd207, 1'b1, 1'b0};
6493: data_out = {8'd11, 8'd207, 1'b1, 1'b0};
6494: data_out = {8'd14, 8'd207, 1'b1, 1'b0};
6495: data_out = {8'd18, 8'd207, 1'b1, 1'b0};
6496: data_out = {8'd21, 8'd207, 1'b1, 1'b0};
6497: data_out = {8'd25, 8'd207, 1'b1, 1'b0};
6498: data_out = {8'd28, 8'd207, 1'b1, 1'b0};
6499: data_out = {8'd32, 8'd207, 1'b1, 1'b0};
6500: data_out = {8'd37, 8'd207, 1'b1, 1'b0};
6501: data_out = {8'd41, 8'd207, 1'b1, 1'b0};
6502: data_out = {8'd45, 8'd207, 1'b1, 1'b0};
6503: data_out = {8'd48, 8'd207, 1'b1, 1'b0};
6504: data_out = {8'd52, 8'd207, 1'b1, 1'b0};
6505: data_out = {8'd61, 8'd207, 1'b1, 1'b0};
6506: data_out = {8'd65, 8'd207, 1'b1, 1'b0};
6507: data_out = {8'd68, 8'd207, 1'b1, 1'b0};
6508: data_out = {8'd72, 8'd207, 1'b1, 1'b0};
6509: data_out = {8'd77, 8'd207, 1'b1, 1'b0};
6510: data_out = {8'd83, 8'd207, 1'b1, 1'b0};
6511: data_out = {8'd87, 8'd207, 1'b1, 1'b0};
6512: data_out = {8'd91, 8'd207, 1'b1, 1'b0};
6513: data_out = {8'd94, 8'd207, 1'b1, 1'b0};
6514: data_out = {8'd98, 8'd207, 1'b1, 1'b0};
6515: data_out = {8'd114, 8'd207, 1'b1, 1'b0};
6516: data_out = {8'd116, 8'd207, 1'b1, 1'b0};
6517: data_out = {8'd119, 8'd207, 1'b1, 1'b0};
6518: data_out = {8'd123, 8'd207, 1'b1, 1'b0};
6519: data_out = {8'd126, 8'd207, 1'b1, 1'b0};
6520: data_out = {8'd130, 8'd207, 1'b1, 1'b0};
6521: data_out = {8'd133, 8'd207, 1'b1, 1'b0};
6522: data_out = {8'd137, 8'd207, 1'b1, 1'b0};
6523: data_out = {8'd141, 8'd207, 1'b1, 1'b0};
6524: data_out = {8'd143, 8'd207, 1'b1, 1'b0};
6525: data_out = {8'd5, 8'd208, 1'b1, 1'b0};
6526: data_out = {8'd8, 8'd208, 1'b1, 1'b0};
6527: data_out = {8'd11, 8'd208, 1'b1, 1'b0};
6528: data_out = {8'd14, 8'd208, 1'b1, 1'b0};
6529: data_out = {8'd18, 8'd208, 1'b1, 1'b0};
6530: data_out = {8'd21, 8'd208, 1'b1, 1'b0};
6531: data_out = {8'd25, 8'd208, 1'b1, 1'b0};
6532: data_out = {8'd28, 8'd208, 1'b1, 1'b0};
6533: data_out = {8'd32, 8'd208, 1'b1, 1'b0};
6534: data_out = {8'd37, 8'd208, 1'b1, 1'b0};
6535: data_out = {8'd41, 8'd208, 1'b1, 1'b0};
6536: data_out = {8'd45, 8'd208, 1'b1, 1'b0};
6537: data_out = {8'd48, 8'd208, 1'b1, 1'b0};
6538: data_out = {8'd61, 8'd208, 1'b1, 1'b0};
6539: data_out = {8'd65, 8'd208, 1'b1, 1'b0};
6540: data_out = {8'd68, 8'd208, 1'b1, 1'b0};
6541: data_out = {8'd72, 8'd208, 1'b1, 1'b0};
6542: data_out = {8'd77, 8'd208, 1'b1, 1'b0};
6543: data_out = {8'd83, 8'd208, 1'b1, 1'b0};
6544: data_out = {8'd87, 8'd208, 1'b1, 1'b0};
6545: data_out = {8'd91, 8'd208, 1'b1, 1'b0};
6546: data_out = {8'd94, 8'd208, 1'b1, 1'b0};
6547: data_out = {8'd98, 8'd208, 1'b1, 1'b0};
6548: data_out = {8'd114, 8'd208, 1'b1, 1'b0};
6549: data_out = {8'd123, 8'd208, 1'b1, 1'b0};
6550: data_out = {8'd126, 8'd208, 1'b1, 1'b0};
6551: data_out = {8'd130, 8'd208, 1'b1, 1'b0};
6552: data_out = {8'd137, 8'd208, 1'b1, 1'b0};
6553: data_out = {8'd141, 8'd208, 1'b1, 1'b0};
6554: data_out = {8'd5, 8'd209, 1'b1, 1'b0};
6555: data_out = {8'd8, 8'd209, 1'b1, 1'b0};
6556: data_out = {8'd11, 8'd209, 1'b1, 1'b0};
6557: data_out = {8'd14, 8'd209, 1'b1, 1'b0};
6558: data_out = {8'd18, 8'd209, 1'b1, 1'b0};
6559: data_out = {8'd21, 8'd209, 1'b1, 1'b0};
6560: data_out = {8'd25, 8'd209, 1'b1, 1'b0};
6561: data_out = {8'd28, 8'd209, 1'b1, 1'b0};
6562: data_out = {8'd32, 8'd209, 1'b1, 1'b0};
6563: data_out = {8'd37, 8'd209, 1'b1, 1'b0};
6564: data_out = {8'd41, 8'd209, 1'b1, 1'b0};
6565: data_out = {8'd42, 8'd209, 1'b1, 1'b0};
6566: data_out = {8'd43, 8'd209, 1'b1, 1'b0};
6567: data_out = {8'd44, 8'd209, 1'b1, 1'b0};
6568: data_out = {8'd48, 8'd209, 1'b1, 1'b0};
6569: data_out = {8'd49, 8'd209, 1'b1, 1'b0};
6570: data_out = {8'd50, 8'd209, 1'b1, 1'b0};
6571: data_out = {8'd51, 8'd209, 1'b1, 1'b0};
6572: data_out = {8'd52, 8'd209, 1'b1, 1'b0};
6573: data_out = {8'd61, 8'd209, 1'b1, 1'b0};
6574: data_out = {8'd65, 8'd209, 1'b1, 1'b0};
6575: data_out = {8'd68, 8'd209, 1'b1, 1'b0};
6576: data_out = {8'd72, 8'd209, 1'b1, 1'b0};
6577: data_out = {8'd77, 8'd209, 1'b1, 1'b0};
6578: data_out = {8'd83, 8'd209, 1'b1, 1'b0};
6579: data_out = {8'd87, 8'd209, 1'b1, 1'b0};
6580: data_out = {8'd91, 8'd209, 1'b1, 1'b0};
6581: data_out = {8'd94, 8'd209, 1'b1, 1'b0};
6582: data_out = {8'd95, 8'd209, 1'b1, 1'b0};
6583: data_out = {8'd96, 8'd209, 1'b1, 1'b0};
6584: data_out = {8'd97, 8'd209, 1'b1, 1'b0};
6585: data_out = {8'd102, 8'd209, 1'b1, 1'b0};
6586: data_out = {8'd114, 8'd209, 1'b1, 1'b0};
6587: data_out = {8'd120, 8'd209, 1'b1, 1'b0};
6588: data_out = {8'd121, 8'd209, 1'b1, 1'b0};
6589: data_out = {8'd122, 8'd209, 1'b1, 1'b0};
6590: data_out = {8'd123, 8'd209, 1'b1, 1'b0};
6591: data_out = {8'd126, 8'd209, 1'b1, 1'b0};
6592: data_out = {8'd130, 8'd209, 1'b1, 1'b0};
6593: data_out = {8'd134, 8'd209, 1'b1, 1'b0};
6594: data_out = {8'd135, 8'd209, 1'b1, 1'b0};
6595: data_out = {8'd136, 8'd209, 1'b1, 1'b0};
6596: data_out = {8'd137, 8'd209, 1'b1, 1'b0};
6597: data_out = {8'd141, 8'd209, 1'b1, 1'b0};
6598: data_out = {8'd148, 8'd209, 1'b1, 1'b0};
6599: data_out = {8'd5, 8'd210, 1'b1, 1'b0};
6600: data_out = {8'd8, 8'd210, 1'b1, 1'b0};
6601: data_out = {8'd11, 8'd210, 1'b1, 1'b0};
6602: data_out = {8'd14, 8'd210, 1'b1, 1'b0};
6603: data_out = {8'd18, 8'd210, 1'b1, 1'b0};
6604: data_out = {8'd21, 8'd210, 1'b1, 1'b0};
6605: data_out = {8'd25, 8'd210, 1'b1, 1'b0};
6606: data_out = {8'd28, 8'd210, 1'b1, 1'b0};
6607: data_out = {8'd32, 8'd210, 1'b1, 1'b0};
6608: data_out = {8'd37, 8'd210, 1'b1, 1'b0};
6609: data_out = {8'd41, 8'd210, 1'b1, 1'b0};
6610: data_out = {8'd52, 8'd210, 1'b1, 1'b0};
6611: data_out = {8'd61, 8'd210, 1'b1, 1'b0};
6612: data_out = {8'd65, 8'd210, 1'b1, 1'b0};
6613: data_out = {8'd68, 8'd210, 1'b1, 1'b0};
6614: data_out = {8'd72, 8'd210, 1'b1, 1'b0};
6615: data_out = {8'd77, 8'd210, 1'b1, 1'b0};
6616: data_out = {8'd83, 8'd210, 1'b1, 1'b0};
6617: data_out = {8'd87, 8'd210, 1'b1, 1'b0};
6618: data_out = {8'd91, 8'd210, 1'b1, 1'b0};
6619: data_out = {8'd94, 8'd210, 1'b1, 1'b0};
6620: data_out = {8'd114, 8'd210, 1'b1, 1'b0};
6621: data_out = {8'd119, 8'd210, 1'b1, 1'b0};
6622: data_out = {8'd123, 8'd210, 1'b1, 1'b0};
6623: data_out = {8'd126, 8'd210, 1'b1, 1'b0};
6624: data_out = {8'd130, 8'd210, 1'b1, 1'b0};
6625: data_out = {8'd133, 8'd210, 1'b1, 1'b0};
6626: data_out = {8'd137, 8'd210, 1'b1, 1'b0};
6627: data_out = {8'd141, 8'd210, 1'b1, 1'b0};
6628: data_out = {8'd5, 8'd211, 1'b1, 1'b0};
6629: data_out = {8'd8, 8'd211, 1'b1, 1'b0};
6630: data_out = {8'd11, 8'd211, 1'b1, 1'b0};
6631: data_out = {8'd14, 8'd211, 1'b1, 1'b0};
6632: data_out = {8'd18, 8'd211, 1'b1, 1'b0};
6633: data_out = {8'd21, 8'd211, 1'b1, 1'b0};
6634: data_out = {8'd25, 8'd211, 1'b1, 1'b0};
6635: data_out = {8'd28, 8'd211, 1'b1, 1'b0};
6636: data_out = {8'd32, 8'd211, 1'b1, 1'b0};
6637: data_out = {8'd37, 8'd211, 1'b1, 1'b0};
6638: data_out = {8'd41, 8'd211, 1'b1, 1'b0};
6639: data_out = {8'd52, 8'd211, 1'b1, 1'b0};
6640: data_out = {8'd61, 8'd211, 1'b1, 1'b0};
6641: data_out = {8'd65, 8'd211, 1'b1, 1'b0};
6642: data_out = {8'd68, 8'd211, 1'b1, 1'b0};
6643: data_out = {8'd72, 8'd211, 1'b1, 1'b0};
6644: data_out = {8'd77, 8'd211, 1'b1, 1'b0};
6645: data_out = {8'd83, 8'd211, 1'b1, 1'b0};
6646: data_out = {8'd87, 8'd211, 1'b1, 1'b0};
6647: data_out = {8'd91, 8'd211, 1'b1, 1'b0};
6648: data_out = {8'd94, 8'd211, 1'b1, 1'b0};
6649: data_out = {8'd114, 8'd211, 1'b1, 1'b0};
6650: data_out = {8'd119, 8'd211, 1'b1, 1'b0};
6651: data_out = {8'd123, 8'd211, 1'b1, 1'b0};
6652: data_out = {8'd126, 8'd211, 1'b1, 1'b0};
6653: data_out = {8'd130, 8'd211, 1'b1, 1'b0};
6654: data_out = {8'd133, 8'd211, 1'b1, 1'b0};
6655: data_out = {8'd137, 8'd211, 1'b1, 1'b0};
6656: data_out = {8'd141, 8'd211, 1'b1, 1'b0};
6657: data_out = {8'd5, 8'd212, 1'b1, 1'b0};
6658: data_out = {8'd8, 8'd212, 1'b1, 1'b0};
6659: data_out = {8'd11, 8'd212, 1'b1, 1'b0};
6660: data_out = {8'd14, 8'd212, 1'b1, 1'b0};
6661: data_out = {8'd15, 8'd212, 1'b1, 1'b0};
6662: data_out = {8'd16, 8'd212, 1'b1, 1'b0};
6663: data_out = {8'd17, 8'd212, 1'b1, 1'b0};
6664: data_out = {8'd18, 8'd212, 1'b1, 1'b0};
6665: data_out = {8'd21, 8'd212, 1'b1, 1'b0};
6666: data_out = {8'd22, 8'd212, 1'b1, 1'b0};
6667: data_out = {8'd23, 8'd212, 1'b1, 1'b0};
6668: data_out = {8'd24, 8'd212, 1'b1, 1'b0};
6669: data_out = {8'd25, 8'd212, 1'b1, 1'b0};
6670: data_out = {8'd28, 8'd212, 1'b1, 1'b0};
6671: data_out = {8'd29, 8'd212, 1'b1, 1'b0};
6672: data_out = {8'd30, 8'd212, 1'b1, 1'b0};
6673: data_out = {8'd31, 8'd212, 1'b1, 1'b0};
6674: data_out = {8'd32, 8'd212, 1'b1, 1'b0};
6675: data_out = {8'd35, 8'd212, 1'b1, 1'b0};
6676: data_out = {8'd36, 8'd212, 1'b1, 1'b0};
6677: data_out = {8'd37, 8'd212, 1'b1, 1'b0};
6678: data_out = {8'd38, 8'd212, 1'b1, 1'b0};
6679: data_out = {8'd39, 8'd212, 1'b1, 1'b0};
6680: data_out = {8'd41, 8'd212, 1'b1, 1'b0};
6681: data_out = {8'd42, 8'd212, 1'b1, 1'b0};
6682: data_out = {8'd43, 8'd212, 1'b1, 1'b0};
6683: data_out = {8'd44, 8'd212, 1'b1, 1'b0};
6684: data_out = {8'd45, 8'd212, 1'b1, 1'b0};
6685: data_out = {8'd48, 8'd212, 1'b1, 1'b0};
6686: data_out = {8'd49, 8'd212, 1'b1, 1'b0};
6687: data_out = {8'd50, 8'd212, 1'b1, 1'b0};
6688: data_out = {8'd51, 8'd212, 1'b1, 1'b0};
6689: data_out = {8'd52, 8'd212, 1'b1, 1'b0};
6690: data_out = {8'd61, 8'd212, 1'b1, 1'b0};
6691: data_out = {8'd62, 8'd212, 1'b1, 1'b0};
6692: data_out = {8'd63, 8'd212, 1'b1, 1'b0};
6693: data_out = {8'd64, 8'd212, 1'b1, 1'b0};
6694: data_out = {8'd65, 8'd212, 1'b1, 1'b0};
6695: data_out = {8'd68, 8'd212, 1'b1, 1'b0};
6696: data_out = {8'd72, 8'd212, 1'b1, 1'b0};
6697: data_out = {8'd75, 8'd212, 1'b1, 1'b0};
6698: data_out = {8'd76, 8'd212, 1'b1, 1'b0};
6699: data_out = {8'd77, 8'd212, 1'b1, 1'b0};
6700: data_out = {8'd78, 8'd212, 1'b1, 1'b0};
6701: data_out = {8'd79, 8'd212, 1'b1, 1'b0};
6702: data_out = {8'd81, 8'd212, 1'b1, 1'b0};
6703: data_out = {8'd82, 8'd212, 1'b1, 1'b0};
6704: data_out = {8'd83, 8'd212, 1'b1, 1'b0};
6705: data_out = {8'd84, 8'd212, 1'b1, 1'b0};
6706: data_out = {8'd85, 8'd212, 1'b1, 1'b0};
6707: data_out = {8'd87, 8'd212, 1'b1, 1'b0};
6708: data_out = {8'd91, 8'd212, 1'b1, 1'b0};
6709: data_out = {8'd94, 8'd212, 1'b1, 1'b0};
6710: data_out = {8'd95, 8'd212, 1'b1, 1'b0};
6711: data_out = {8'd96, 8'd212, 1'b1, 1'b0};
6712: data_out = {8'd97, 8'd212, 1'b1, 1'b0};
6713: data_out = {8'd98, 8'd212, 1'b1, 1'b0};
6714: data_out = {8'd102, 8'd212, 1'b1, 1'b0};
6715: data_out = {8'd112, 8'd212, 1'b1, 1'b0};
6716: data_out = {8'd113, 8'd212, 1'b1, 1'b0};
6717: data_out = {8'd114, 8'd212, 1'b1, 1'b0};
6718: data_out = {8'd115, 8'd212, 1'b1, 1'b0};
6719: data_out = {8'd116, 8'd212, 1'b1, 1'b0};
6720: data_out = {8'd117, 8'd212, 1'b1, 1'b0};
6721: data_out = {8'd119, 8'd212, 1'b1, 1'b0};
6722: data_out = {8'd120, 8'd212, 1'b1, 1'b0};
6723: data_out = {8'd121, 8'd212, 1'b1, 1'b0};
6724: data_out = {8'd122, 8'd212, 1'b1, 1'b0};
6725: data_out = {8'd123, 8'd212, 1'b1, 1'b0};
6726: data_out = {8'd126, 8'd212, 1'b1, 1'b0};
6727: data_out = {8'd127, 8'd212, 1'b1, 1'b0};
6728: data_out = {8'd128, 8'd212, 1'b1, 1'b0};
6729: data_out = {8'd129, 8'd212, 1'b1, 1'b0};
6730: data_out = {8'd130, 8'd212, 1'b1, 1'b0};
6731: data_out = {8'd133, 8'd212, 1'b1, 1'b0};
6732: data_out = {8'd134, 8'd212, 1'b1, 1'b0};
6733: data_out = {8'd135, 8'd212, 1'b1, 1'b0};
6734: data_out = {8'd136, 8'd212, 1'b1, 1'b0};
6735: data_out = {8'd137, 8'd212, 1'b1, 1'b0};
6736: data_out = {8'd139, 8'd212, 1'b1, 1'b0};
6737: data_out = {8'd140, 8'd212, 1'b1, 1'b0};
6738: data_out = {8'd141, 8'd212, 1'b1, 1'b0};
6739: data_out = {8'd142, 8'd212, 1'b1, 1'b0};
6740: data_out = {8'd143, 8'd212, 1'b1, 1'b0};
6741: data_out = {8'd144, 8'd212, 1'b1, 1'b0};
6742: data_out = {8'd148, 8'd212, 1'b1, 1'b0};
6743: data_out = {8'd147, 8'd213, 1'b1, 1'b0};
6744: data_out = {8'd148, 8'd213, 1'b1, 1'b0};
6745: data_out = {8'd124, 8'd217, 1'b1, 1'b0};
6746: data_out = {8'd144, 8'd217, 1'b1, 1'b0};
6747: data_out = {8'd148, 8'd217, 1'b1, 1'b0};
6748: data_out = {8'd149, 8'd217, 1'b1, 1'b0};
6749: data_out = {8'd150, 8'd217, 1'b1, 1'b0};
6750: data_out = {8'd183, 8'd217, 1'b1, 1'b0};
6751: data_out = {8'd191, 8'd217, 1'b1, 1'b0};
6752: data_out = {8'd150, 8'd218, 1'b1, 1'b0};
6753: data_out = {8'd191, 8'd218, 1'b1, 1'b0};
6754: data_out = {8'd113, 8'd219, 1'b1, 1'b0};
6755: data_out = {8'd114, 8'd219, 1'b1, 1'b0};
6756: data_out = {8'd115, 8'd219, 1'b1, 1'b0};
6757: data_out = {8'd116, 8'd219, 1'b1, 1'b0};
6758: data_out = {8'd117, 8'd219, 1'b1, 1'b0};
6759: data_out = {8'd118, 8'd219, 1'b1, 1'b0};
6760: data_out = {8'd119, 8'd219, 1'b1, 1'b0};
6761: data_out = {8'd122, 8'd219, 1'b1, 1'b0};
6762: data_out = {8'd123, 8'd219, 1'b1, 1'b0};
6763: data_out = {8'd124, 8'd219, 1'b1, 1'b0};
6764: data_out = {8'd128, 8'd219, 1'b1, 1'b0};
6765: data_out = {8'd129, 8'd219, 1'b1, 1'b0};
6766: data_out = {8'd130, 8'd219, 1'b1, 1'b0};
6767: data_out = {8'd131, 8'd219, 1'b1, 1'b0};
6768: data_out = {8'd132, 8'd219, 1'b1, 1'b0};
6769: data_out = {8'd135, 8'd219, 1'b1, 1'b0};
6770: data_out = {8'd136, 8'd219, 1'b1, 1'b0};
6771: data_out = {8'd137, 8'd219, 1'b1, 1'b0};
6772: data_out = {8'd138, 8'd219, 1'b1, 1'b0};
6773: data_out = {8'd139, 8'd219, 1'b1, 1'b0};
6774: data_out = {8'd142, 8'd219, 1'b1, 1'b0};
6775: data_out = {8'd143, 8'd219, 1'b1, 1'b0};
6776: data_out = {8'd144, 8'd219, 1'b1, 1'b0};
6777: data_out = {8'd150, 8'd219, 1'b1, 1'b0};
6778: data_out = {8'd154, 8'd219, 1'b1, 1'b0};
6779: data_out = {8'd155, 8'd219, 1'b1, 1'b0};
6780: data_out = {8'd156, 8'd219, 1'b1, 1'b0};
6781: data_out = {8'd157, 8'd219, 1'b1, 1'b0};
6782: data_out = {8'd158, 8'd219, 1'b1, 1'b0};
6783: data_out = {8'd167, 8'd219, 1'b1, 1'b0};
6784: data_out = {8'd168, 8'd219, 1'b1, 1'b0};
6785: data_out = {8'd169, 8'd219, 1'b1, 1'b0};
6786: data_out = {8'd170, 8'd219, 1'b1, 1'b0};
6787: data_out = {8'd171, 8'd219, 1'b1, 1'b0};
6788: data_out = {8'd174, 8'd219, 1'b1, 1'b0};
6789: data_out = {8'd178, 8'd219, 1'b1, 1'b0};
6790: data_out = {8'd181, 8'd219, 1'b1, 1'b0};
6791: data_out = {8'd182, 8'd219, 1'b1, 1'b0};
6792: data_out = {8'd183, 8'd219, 1'b1, 1'b0};
6793: data_out = {8'd187, 8'd219, 1'b1, 1'b0};
6794: data_out = {8'd188, 8'd219, 1'b1, 1'b0};
6795: data_out = {8'd189, 8'd219, 1'b1, 1'b0};
6796: data_out = {8'd190, 8'd219, 1'b1, 1'b0};
6797: data_out = {8'd191, 8'd219, 1'b1, 1'b0};
6798: data_out = {8'd194, 8'd219, 1'b1, 1'b0};
6799: data_out = {8'd195, 8'd219, 1'b1, 1'b0};
6800: data_out = {8'd196, 8'd219, 1'b1, 1'b0};
6801: data_out = {8'd197, 8'd219, 1'b1, 1'b0};
6802: data_out = {8'd198, 8'd219, 1'b1, 1'b0};
6803: data_out = {8'd201, 8'd219, 1'b1, 1'b0};
6804: data_out = {8'd202, 8'd219, 1'b1, 1'b0};
6805: data_out = {8'd203, 8'd219, 1'b1, 1'b0};
6806: data_out = {8'd204, 8'd219, 1'b1, 1'b0};
6807: data_out = {8'd205, 8'd219, 1'b1, 1'b0};
6808: data_out = {8'd208, 8'd219, 1'b1, 1'b0};
6809: data_out = {8'd209, 8'd219, 1'b1, 1'b0};
6810: data_out = {8'd210, 8'd219, 1'b1, 1'b0};
6811: data_out = {8'd211, 8'd219, 1'b1, 1'b0};
6812: data_out = {8'd212, 8'd219, 1'b1, 1'b0};
6813: data_out = {8'd215, 8'd219, 1'b1, 1'b0};
6814: data_out = {8'd216, 8'd219, 1'b1, 1'b0};
6815: data_out = {8'd217, 8'd219, 1'b1, 1'b0};
6816: data_out = {8'd218, 8'd219, 1'b1, 1'b0};
6817: data_out = {8'd219, 8'd219, 1'b1, 1'b0};
6818: data_out = {8'd113, 8'd220, 1'b1, 1'b0};
6819: data_out = {8'd116, 8'd220, 1'b1, 1'b0};
6820: data_out = {8'd119, 8'd220, 1'b1, 1'b0};
6821: data_out = {8'd124, 8'd220, 1'b1, 1'b0};
6822: data_out = {8'd128, 8'd220, 1'b1, 1'b0};
6823: data_out = {8'd132, 8'd220, 1'b1, 1'b0};
6824: data_out = {8'd135, 8'd220, 1'b1, 1'b0};
6825: data_out = {8'd139, 8'd220, 1'b1, 1'b0};
6826: data_out = {8'd144, 8'd220, 1'b1, 1'b0};
6827: data_out = {8'd150, 8'd220, 1'b1, 1'b0};
6828: data_out = {8'd154, 8'd220, 1'b1, 1'b0};
6829: data_out = {8'd158, 8'd220, 1'b1, 1'b0};
6830: data_out = {8'd167, 8'd220, 1'b1, 1'b0};
6831: data_out = {8'd170, 8'd220, 1'b1, 1'b0};
6832: data_out = {8'd174, 8'd220, 1'b1, 1'b0};
6833: data_out = {8'd178, 8'd220, 1'b1, 1'b0};
6834: data_out = {8'd183, 8'd220, 1'b1, 1'b0};
6835: data_out = {8'd187, 8'd220, 1'b1, 1'b0};
6836: data_out = {8'd191, 8'd220, 1'b1, 1'b0};
6837: data_out = {8'd194, 8'd220, 1'b1, 1'b0};
6838: data_out = {8'd198, 8'd220, 1'b1, 1'b0};
6839: data_out = {8'd201, 8'd220, 1'b1, 1'b0};
6840: data_out = {8'd205, 8'd220, 1'b1, 1'b0};
6841: data_out = {8'd208, 8'd220, 1'b1, 1'b0};
6842: data_out = {8'd212, 8'd220, 1'b1, 1'b0};
6843: data_out = {8'd215, 8'd220, 1'b1, 1'b0};
6844: data_out = {8'd219, 8'd220, 1'b1, 1'b0};
6845: data_out = {8'd113, 8'd221, 1'b1, 1'b0};
6846: data_out = {8'd116, 8'd221, 1'b1, 1'b0};
6847: data_out = {8'd119, 8'd221, 1'b1, 1'b0};
6848: data_out = {8'd124, 8'd221, 1'b1, 1'b0};
6849: data_out = {8'd128, 8'd221, 1'b1, 1'b0};
6850: data_out = {8'd135, 8'd221, 1'b1, 1'b0};
6851: data_out = {8'd144, 8'd221, 1'b1, 1'b0};
6852: data_out = {8'd150, 8'd221, 1'b1, 1'b0};
6853: data_out = {8'd154, 8'd221, 1'b1, 1'b0};
6854: data_out = {8'd158, 8'd221, 1'b1, 1'b0};
6855: data_out = {8'd167, 8'd221, 1'b1, 1'b0};
6856: data_out = {8'd170, 8'd221, 1'b1, 1'b0};
6857: data_out = {8'd174, 8'd221, 1'b1, 1'b0};
6858: data_out = {8'd178, 8'd221, 1'b1, 1'b0};
6859: data_out = {8'd183, 8'd221, 1'b1, 1'b0};
6860: data_out = {8'd187, 8'd221, 1'b1, 1'b0};
6861: data_out = {8'd191, 8'd221, 1'b1, 1'b0};
6862: data_out = {8'd198, 8'd221, 1'b1, 1'b0};
6863: data_out = {8'd201, 8'd221, 1'b1, 1'b0};
6864: data_out = {8'd205, 8'd221, 1'b1, 1'b0};
6865: data_out = {8'd208, 8'd221, 1'b1, 1'b0};
6866: data_out = {8'd215, 8'd221, 1'b1, 1'b0};
6867: data_out = {8'd219, 8'd221, 1'b1, 1'b0};
6868: data_out = {8'd113, 8'd222, 1'b1, 1'b0};
6869: data_out = {8'd116, 8'd222, 1'b1, 1'b0};
6870: data_out = {8'd119, 8'd222, 1'b1, 1'b0};
6871: data_out = {8'd124, 8'd222, 1'b1, 1'b0};
6872: data_out = {8'd128, 8'd222, 1'b1, 1'b0};
6873: data_out = {8'd129, 8'd222, 1'b1, 1'b0};
6874: data_out = {8'd130, 8'd222, 1'b1, 1'b0};
6875: data_out = {8'd131, 8'd222, 1'b1, 1'b0};
6876: data_out = {8'd132, 8'd222, 1'b1, 1'b0};
6877: data_out = {8'd135, 8'd222, 1'b1, 1'b0};
6878: data_out = {8'd136, 8'd222, 1'b1, 1'b0};
6879: data_out = {8'd137, 8'd222, 1'b1, 1'b0};
6880: data_out = {8'd138, 8'd222, 1'b1, 1'b0};
6881: data_out = {8'd139, 8'd222, 1'b1, 1'b0};
6882: data_out = {8'd144, 8'd222, 1'b1, 1'b0};
6883: data_out = {8'd150, 8'd222, 1'b1, 1'b0};
6884: data_out = {8'd154, 8'd222, 1'b1, 1'b0};
6885: data_out = {8'd155, 8'd222, 1'b1, 1'b0};
6886: data_out = {8'd156, 8'd222, 1'b1, 1'b0};
6887: data_out = {8'd157, 8'd222, 1'b1, 1'b0};
6888: data_out = {8'd167, 8'd222, 1'b1, 1'b0};
6889: data_out = {8'd170, 8'd222, 1'b1, 1'b0};
6890: data_out = {8'd174, 8'd222, 1'b1, 1'b0};
6891: data_out = {8'd178, 8'd222, 1'b1, 1'b0};
6892: data_out = {8'd183, 8'd222, 1'b1, 1'b0};
6893: data_out = {8'd187, 8'd222, 1'b1, 1'b0};
6894: data_out = {8'd191, 8'd222, 1'b1, 1'b0};
6895: data_out = {8'd195, 8'd222, 1'b1, 1'b0};
6896: data_out = {8'd196, 8'd222, 1'b1, 1'b0};
6897: data_out = {8'd197, 8'd222, 1'b1, 1'b0};
6898: data_out = {8'd198, 8'd222, 1'b1, 1'b0};
6899: data_out = {8'd201, 8'd222, 1'b1, 1'b0};
6900: data_out = {8'd205, 8'd222, 1'b1, 1'b0};
6901: data_out = {8'd208, 8'd222, 1'b1, 1'b0};
6902: data_out = {8'd215, 8'd222, 1'b1, 1'b0};
6903: data_out = {8'd216, 8'd222, 1'b1, 1'b0};
6904: data_out = {8'd217, 8'd222, 1'b1, 1'b0};
6905: data_out = {8'd218, 8'd222, 1'b1, 1'b0};
6906: data_out = {8'd224, 8'd222, 1'b1, 1'b0};
6907: data_out = {8'd113, 8'd223, 1'b1, 1'b0};
6908: data_out = {8'd116, 8'd223, 1'b1, 1'b0};
6909: data_out = {8'd119, 8'd223, 1'b1, 1'b0};
6910: data_out = {8'd124, 8'd223, 1'b1, 1'b0};
6911: data_out = {8'd132, 8'd223, 1'b1, 1'b0};
6912: data_out = {8'd139, 8'd223, 1'b1, 1'b0};
6913: data_out = {8'd144, 8'd223, 1'b1, 1'b0};
6914: data_out = {8'd150, 8'd223, 1'b1, 1'b0};
6915: data_out = {8'd154, 8'd223, 1'b1, 1'b0};
6916: data_out = {8'd167, 8'd223, 1'b1, 1'b0};
6917: data_out = {8'd168, 8'd223, 1'b1, 1'b0};
6918: data_out = {8'd169, 8'd223, 1'b1, 1'b0};
6919: data_out = {8'd170, 8'd223, 1'b1, 1'b0};
6920: data_out = {8'd174, 8'd223, 1'b1, 1'b0};
6921: data_out = {8'd178, 8'd223, 1'b1, 1'b0};
6922: data_out = {8'd183, 8'd223, 1'b1, 1'b0};
6923: data_out = {8'd187, 8'd223, 1'b1, 1'b0};
6924: data_out = {8'd191, 8'd223, 1'b1, 1'b0};
6925: data_out = {8'd194, 8'd223, 1'b1, 1'b0};
6926: data_out = {8'd198, 8'd223, 1'b1, 1'b0};
6927: data_out = {8'd201, 8'd223, 1'b1, 1'b0};
6928: data_out = {8'd205, 8'd223, 1'b1, 1'b0};
6929: data_out = {8'd208, 8'd223, 1'b1, 1'b0};
6930: data_out = {8'd215, 8'd223, 1'b1, 1'b0};
6931: data_out = {8'd113, 8'd224, 1'b1, 1'b0};
6932: data_out = {8'd116, 8'd224, 1'b1, 1'b0};
6933: data_out = {8'd119, 8'd224, 1'b1, 1'b0};
6934: data_out = {8'd124, 8'd224, 1'b1, 1'b0};
6935: data_out = {8'd132, 8'd224, 1'b1, 1'b0};
6936: data_out = {8'd139, 8'd224, 1'b1, 1'b0};
6937: data_out = {8'd144, 8'd224, 1'b1, 1'b0};
6938: data_out = {8'd150, 8'd224, 1'b1, 1'b0};
6939: data_out = {8'd154, 8'd224, 1'b1, 1'b0};
6940: data_out = {8'd167, 8'd224, 1'b1, 1'b0};
6941: data_out = {8'd174, 8'd224, 1'b1, 1'b0};
6942: data_out = {8'd178, 8'd224, 1'b1, 1'b0};
6943: data_out = {8'd183, 8'd224, 1'b1, 1'b0};
6944: data_out = {8'd187, 8'd224, 1'b1, 1'b0};
6945: data_out = {8'd191, 8'd224, 1'b1, 1'b0};
6946: data_out = {8'd194, 8'd224, 1'b1, 1'b0};
6947: data_out = {8'd198, 8'd224, 1'b1, 1'b0};
6948: data_out = {8'd201, 8'd224, 1'b1, 1'b0};
6949: data_out = {8'd205, 8'd224, 1'b1, 1'b0};
6950: data_out = {8'd208, 8'd224, 1'b1, 1'b0};
6951: data_out = {8'd215, 8'd224, 1'b1, 1'b0};
6952: data_out = {8'd113, 8'd225, 1'b1, 1'b0};
6953: data_out = {8'd116, 8'd225, 1'b1, 1'b0};
6954: data_out = {8'd119, 8'd225, 1'b1, 1'b0};
6955: data_out = {8'd122, 8'd225, 1'b1, 1'b0};
6956: data_out = {8'd123, 8'd225, 1'b1, 1'b0};
6957: data_out = {8'd124, 8'd225, 1'b1, 1'b0};
6958: data_out = {8'd125, 8'd225, 1'b1, 1'b0};
6959: data_out = {8'd126, 8'd225, 1'b1, 1'b0};
6960: data_out = {8'd128, 8'd225, 1'b1, 1'b0};
6961: data_out = {8'd129, 8'd225, 1'b1, 1'b0};
6962: data_out = {8'd130, 8'd225, 1'b1, 1'b0};
6963: data_out = {8'd131, 8'd225, 1'b1, 1'b0};
6964: data_out = {8'd132, 8'd225, 1'b1, 1'b0};
6965: data_out = {8'd135, 8'd225, 1'b1, 1'b0};
6966: data_out = {8'd136, 8'd225, 1'b1, 1'b0};
6967: data_out = {8'd137, 8'd225, 1'b1, 1'b0};
6968: data_out = {8'd138, 8'd225, 1'b1, 1'b0};
6969: data_out = {8'd139, 8'd225, 1'b1, 1'b0};
6970: data_out = {8'd142, 8'd225, 1'b1, 1'b0};
6971: data_out = {8'd143, 8'd225, 1'b1, 1'b0};
6972: data_out = {8'd144, 8'd225, 1'b1, 1'b0};
6973: data_out = {8'd145, 8'd225, 1'b1, 1'b0};
6974: data_out = {8'd146, 8'd225, 1'b1, 1'b0};
6975: data_out = {8'd148, 8'd225, 1'b1, 1'b0};
6976: data_out = {8'd149, 8'd225, 1'b1, 1'b0};
6977: data_out = {8'd150, 8'd225, 1'b1, 1'b0};
6978: data_out = {8'd151, 8'd225, 1'b1, 1'b0};
6979: data_out = {8'd152, 8'd225, 1'b1, 1'b0};
6980: data_out = {8'd154, 8'd225, 1'b1, 1'b0};
6981: data_out = {8'd155, 8'd225, 1'b1, 1'b0};
6982: data_out = {8'd156, 8'd225, 1'b1, 1'b0};
6983: data_out = {8'd157, 8'd225, 1'b1, 1'b0};
6984: data_out = {8'd158, 8'd225, 1'b1, 1'b0};
6985: data_out = {8'd167, 8'd225, 1'b1, 1'b0};
6986: data_out = {8'd168, 8'd225, 1'b1, 1'b0};
6987: data_out = {8'd169, 8'd225, 1'b1, 1'b0};
6988: data_out = {8'd170, 8'd225, 1'b1, 1'b0};
6989: data_out = {8'd171, 8'd225, 1'b1, 1'b0};
6990: data_out = {8'd174, 8'd225, 1'b1, 1'b0};
6991: data_out = {8'd175, 8'd225, 1'b1, 1'b0};
6992: data_out = {8'd176, 8'd225, 1'b1, 1'b0};
6993: data_out = {8'd177, 8'd225, 1'b1, 1'b0};
6994: data_out = {8'd178, 8'd225, 1'b1, 1'b0};
6995: data_out = {8'd181, 8'd225, 1'b1, 1'b0};
6996: data_out = {8'd182, 8'd225, 1'b1, 1'b0};
6997: data_out = {8'd183, 8'd225, 1'b1, 1'b0};
6998: data_out = {8'd184, 8'd225, 1'b1, 1'b0};
6999: data_out = {8'd185, 8'd225, 1'b1, 1'b0};
7000: data_out = {8'd187, 8'd225, 1'b1, 1'b0};
7001: data_out = {8'd188, 8'd225, 1'b1, 1'b0};
7002: data_out = {8'd189, 8'd225, 1'b1, 1'b0};
7003: data_out = {8'd190, 8'd225, 1'b1, 1'b0};
7004: data_out = {8'd191, 8'd225, 1'b1, 1'b0};
7005: data_out = {8'd194, 8'd225, 1'b1, 1'b0};
7006: data_out = {8'd195, 8'd225, 1'b1, 1'b0};
7007: data_out = {8'd196, 8'd225, 1'b1, 1'b0};
7008: data_out = {8'd197, 8'd225, 1'b1, 1'b0};
7009: data_out = {8'd198, 8'd225, 1'b1, 1'b0};
7010: data_out = {8'd201, 8'd225, 1'b1, 1'b0};
7011: data_out = {8'd205, 8'd225, 1'b1, 1'b0};
7012: data_out = {8'd208, 8'd225, 1'b1, 1'b0};
7013: data_out = {8'd209, 8'd225, 1'b1, 1'b0};
7014: data_out = {8'd210, 8'd225, 1'b1, 1'b0};
7015: data_out = {8'd211, 8'd225, 1'b1, 1'b0};
7016: data_out = {8'd212, 8'd225, 1'b1, 1'b0};
7017: data_out = {8'd215, 8'd225, 1'b1, 1'b0};
7018: data_out = {8'd216, 8'd225, 1'b1, 1'b0};
7019: data_out = {8'd217, 8'd225, 1'b1, 1'b0};
7020: data_out = {8'd218, 8'd225, 1'b1, 1'b0};
7021: data_out = {8'd219, 8'd225, 1'b1, 1'b0};
7022: data_out = {8'd224, 8'd225, 1'b1, 1'b0};
7023: data_out = {8'd167, 8'd226, 1'b1, 1'b0};
7024: data_out = {8'd171, 8'd226, 1'b1, 1'b0};
7025: data_out = {8'd223, 8'd226, 1'b1, 1'b0};
7026: data_out = {8'd224, 8'd226, 1'b1, 1'b0};
7027: data_out = {8'd167, 8'd227, 1'b1, 1'b0};
7028: data_out = {8'd171, 8'd227, 1'b1, 1'b0};
7029: data_out = {8'd167, 8'd228, 1'b1, 1'b0};
7030: data_out = {8'd168, 8'd228, 1'b1, 1'b0};
7031: data_out = {8'd169, 8'd228, 1'b1, 1'b0};
7032: data_out = {8'd170, 8'd228, 1'b1, 1'b0};
7033: data_out = {8'd171, 8'd228, 1'b1, 1'b0};
7034: data_out = {8'd217, 8'd243, 1'b1, 1'b0};
7035: data_out = {8'd226, 8'd243, 1'b1, 1'b0};
7036: data_out = {8'd227, 8'd243, 1'b1, 1'b0};
7037: data_out = {8'd228, 8'd243, 1'b1, 1'b0};
7038: data_out = {8'd246, 8'd243, 1'b1, 1'b0};
7039: data_out = {8'd217, 8'd244, 1'b1, 1'b0};
7040: data_out = {8'd228, 8'd244, 1'b1, 1'b0};
7041: data_out = {8'd246, 8'd244, 1'b1, 1'b0};
7042: data_out = {8'd192, 8'd245, 1'b1, 1'b0};
7043: data_out = {8'd193, 8'd245, 1'b1, 1'b0};
7044: data_out = {8'd194, 8'd245, 1'b1, 1'b0};
7045: data_out = {8'd195, 8'd245, 1'b1, 1'b0};
7046: data_out = {8'd196, 8'd245, 1'b1, 1'b0};
7047: data_out = {8'd199, 8'd245, 1'b1, 1'b0};
7048: data_out = {8'd200, 8'd245, 1'b1, 1'b0};
7049: data_out = {8'd201, 8'd245, 1'b1, 1'b0};
7050: data_out = {8'd202, 8'd245, 1'b1, 1'b0};
7051: data_out = {8'd203, 8'd245, 1'b1, 1'b0};
7052: data_out = {8'd206, 8'd245, 1'b1, 1'b0};
7053: data_out = {8'd207, 8'd245, 1'b1, 1'b0};
7054: data_out = {8'd208, 8'd245, 1'b1, 1'b0};
7055: data_out = {8'd209, 8'd245, 1'b1, 1'b0};
7056: data_out = {8'd210, 8'd245, 1'b1, 1'b0};
7057: data_out = {8'd213, 8'd245, 1'b1, 1'b0};
7058: data_out = {8'd214, 8'd245, 1'b1, 1'b0};
7059: data_out = {8'd215, 8'd245, 1'b1, 1'b0};
7060: data_out = {8'd216, 8'd245, 1'b1, 1'b0};
7061: data_out = {8'd217, 8'd245, 1'b1, 1'b0};
7062: data_out = {8'd228, 8'd245, 1'b1, 1'b0};
7063: data_out = {8'd232, 8'd245, 1'b1, 1'b0};
7064: data_out = {8'd236, 8'd245, 1'b1, 1'b0};
7065: data_out = {8'd239, 8'd245, 1'b1, 1'b0};
7066: data_out = {8'd240, 8'd245, 1'b1, 1'b0};
7067: data_out = {8'd241, 8'd245, 1'b1, 1'b0};
7068: data_out = {8'd242, 8'd245, 1'b1, 1'b0};
7069: data_out = {8'd243, 8'd245, 1'b1, 1'b0};
7070: data_out = {8'd246, 8'd245, 1'b1, 1'b0};
7071: data_out = {8'd250, 8'd245, 1'b1, 1'b0};
7072: data_out = {8'd192, 8'd246, 1'b1, 1'b0};
7073: data_out = {8'd195, 8'd246, 1'b1, 1'b0};
7074: data_out = {8'd199, 8'd246, 1'b1, 1'b0};
7075: data_out = {8'd203, 8'd246, 1'b1, 1'b0};
7076: data_out = {8'd206, 8'd246, 1'b1, 1'b0};
7077: data_out = {8'd210, 8'd246, 1'b1, 1'b0};
7078: data_out = {8'd213, 8'd246, 1'b1, 1'b0};
7079: data_out = {8'd217, 8'd246, 1'b1, 1'b0};
7080: data_out = {8'd228, 8'd246, 1'b1, 1'b0};
7081: data_out = {8'd232, 8'd246, 1'b1, 1'b0};
7082: data_out = {8'd236, 8'd246, 1'b1, 1'b0};
7083: data_out = {8'd239, 8'd246, 1'b1, 1'b0};
7084: data_out = {8'd243, 8'd246, 1'b1, 1'b0};
7085: data_out = {8'd246, 8'd246, 1'b1, 1'b0};
7086: data_out = {8'd249, 8'd246, 1'b1, 1'b0};
7087: data_out = {8'd250, 8'd246, 1'b1, 1'b0};
7088: data_out = {8'd192, 8'd247, 1'b1, 1'b0};
7089: data_out = {8'd195, 8'd247, 1'b1, 1'b0};
7090: data_out = {8'd199, 8'd247, 1'b1, 1'b0};
7091: data_out = {8'd203, 8'd247, 1'b1, 1'b0};
7092: data_out = {8'd206, 8'd247, 1'b1, 1'b0};
7093: data_out = {8'd210, 8'd247, 1'b1, 1'b0};
7094: data_out = {8'd213, 8'd247, 1'b1, 1'b0};
7095: data_out = {8'd217, 8'd247, 1'b1, 1'b0};
7096: data_out = {8'd228, 8'd247, 1'b1, 1'b0};
7097: data_out = {8'd232, 8'd247, 1'b1, 1'b0};
7098: data_out = {8'd236, 8'd247, 1'b1, 1'b0};
7099: data_out = {8'd239, 8'd247, 1'b1, 1'b0};
7100: data_out = {8'd246, 8'd247, 1'b1, 1'b0};
7101: data_out = {8'd249, 8'd247, 1'b1, 1'b0};
7102: data_out = {8'd192, 8'd248, 1'b1, 1'b0};
7103: data_out = {8'd195, 8'd248, 1'b1, 1'b0};
7104: data_out = {8'd199, 8'd248, 1'b1, 1'b0};
7105: data_out = {8'd203, 8'd248, 1'b1, 1'b0};
7106: data_out = {8'd206, 8'd248, 1'b1, 1'b0};
7107: data_out = {8'd210, 8'd248, 1'b1, 1'b0};
7108: data_out = {8'd213, 8'd248, 1'b1, 1'b0};
7109: data_out = {8'd217, 8'd248, 1'b1, 1'b0};
7110: data_out = {8'd228, 8'd248, 1'b1, 1'b0};
7111: data_out = {8'd232, 8'd248, 1'b1, 1'b0};
7112: data_out = {8'd236, 8'd248, 1'b1, 1'b0};
7113: data_out = {8'd239, 8'd248, 1'b1, 1'b0};
7114: data_out = {8'd246, 8'd248, 1'b1, 1'b0};
7115: data_out = {8'd247, 8'd248, 1'b1, 1'b0};
7116: data_out = {8'd248, 8'd248, 1'b1, 1'b0};
7117: data_out = {8'd192, 8'd249, 1'b1, 1'b0};
7118: data_out = {8'd193, 8'd249, 1'b1, 1'b0};
7119: data_out = {8'd194, 8'd249, 1'b1, 1'b0};
7120: data_out = {8'd195, 8'd249, 1'b1, 1'b0};
7121: data_out = {8'd199, 8'd249, 1'b1, 1'b0};
7122: data_out = {8'd203, 8'd249, 1'b1, 1'b0};
7123: data_out = {8'd206, 8'd249, 1'b1, 1'b0};
7124: data_out = {8'd210, 8'd249, 1'b1, 1'b0};
7125: data_out = {8'd213, 8'd249, 1'b1, 1'b0};
7126: data_out = {8'd217, 8'd249, 1'b1, 1'b0};
7127: data_out = {8'd228, 8'd249, 1'b1, 1'b0};
7128: data_out = {8'd232, 8'd249, 1'b1, 1'b0};
7129: data_out = {8'd236, 8'd249, 1'b1, 1'b0};
7130: data_out = {8'd239, 8'd249, 1'b1, 1'b0};
7131: data_out = {8'd246, 8'd249, 1'b1, 1'b0};
7132: data_out = {8'd249, 8'd249, 1'b1, 1'b0};
7133: data_out = {8'd192, 8'd250, 1'b1, 1'b0};
7134: data_out = {8'd199, 8'd250, 1'b1, 1'b0};
7135: data_out = {8'd203, 8'd250, 1'b1, 1'b0};
7136: data_out = {8'd206, 8'd250, 1'b1, 1'b0};
7137: data_out = {8'd210, 8'd250, 1'b1, 1'b0};
7138: data_out = {8'd213, 8'd250, 1'b1, 1'b0};
7139: data_out = {8'd217, 8'd250, 1'b1, 1'b0};
7140: data_out = {8'd228, 8'd250, 1'b1, 1'b0};
7141: data_out = {8'd232, 8'd250, 1'b1, 1'b0};
7142: data_out = {8'd236, 8'd250, 1'b1, 1'b0};
7143: data_out = {8'd239, 8'd250, 1'b1, 1'b0};
7144: data_out = {8'd246, 8'd250, 1'b1, 1'b0};
7145: data_out = {8'd249, 8'd250, 1'b1, 1'b0};
7146: data_out = {8'd250, 8'd250, 1'b1, 1'b0};
7147: data_out = {8'd192, 8'd251, 1'b1, 1'b0};
7148: data_out = {8'd193, 8'd251, 1'b1, 1'b0};
7149: data_out = {8'd194, 8'd251, 1'b1, 1'b0};
7150: data_out = {8'd195, 8'd251, 1'b1, 1'b0};
7151: data_out = {8'd196, 8'd251, 1'b1, 1'b0};
7152: data_out = {8'd199, 8'd251, 1'b1, 1'b0};
7153: data_out = {8'd200, 8'd251, 1'b1, 1'b0};
7154: data_out = {8'd201, 8'd251, 1'b1, 1'b0};
7155: data_out = {8'd202, 8'd251, 1'b1, 1'b0};
7156: data_out = {8'd203, 8'd251, 1'b1, 1'b0};
7157: data_out = {8'd206, 8'd251, 1'b1, 1'b0};
7158: data_out = {8'd207, 8'd251, 1'b1, 1'b0};
7159: data_out = {8'd208, 8'd251, 1'b1, 1'b0};
7160: data_out = {8'd209, 8'd251, 1'b1, 1'b0};
7161: data_out = {8'd210, 8'd251, 1'b1, 1'b0};
7162: data_out = {8'd213, 8'd251, 1'b1, 1'b0};
7163: data_out = {8'd214, 8'd251, 1'b1, 1'b0};
7164: data_out = {8'd215, 8'd251, 1'b1, 1'b0};
7165: data_out = {8'd216, 8'd251, 1'b1, 1'b0};
7166: data_out = {8'd217, 8'd251, 1'b1, 1'b0};
7167: data_out = {8'd226, 8'd251, 1'b1, 1'b0};
7168: data_out = {8'd227, 8'd251, 1'b1, 1'b0};
7169: data_out = {8'd228, 8'd251, 1'b1, 1'b0};
7170: data_out = {8'd229, 8'd251, 1'b1, 1'b0};
7171: data_out = {8'd230, 8'd251, 1'b1, 1'b0};
7172: data_out = {8'd232, 8'd251, 1'b1, 1'b0};
7173: data_out = {8'd233, 8'd251, 1'b1, 1'b0};
7174: data_out = {8'd234, 8'd251, 1'b1, 1'b0};
7175: data_out = {8'd235, 8'd251, 1'b1, 1'b0};
7176: data_out = {8'd236, 8'd251, 1'b1, 1'b0};
7177: data_out = {8'd239, 8'd251, 1'b1, 1'b0};
7178: data_out = {8'd240, 8'd251, 1'b1, 1'b0};
7179: data_out = {8'd241, 8'd251, 1'b1, 1'b0};
7180: data_out = {8'd242, 8'd251, 1'b1, 1'b0};
7181: data_out = {8'd243, 8'd251, 1'b1, 1'b0};
7182: data_out = {8'd246, 8'd251, 1'b1, 1'b0};
7183: data_out = {8'd250, 8'd251, 1'b1, 1'b0};
7184: data_out = {8'd192, 8'd252, 1'b1, 1'b0};
7185: data_out = {8'd196, 8'd252, 1'b1, 1'b0};
7186: data_out = {8'd192, 8'd253, 1'b1, 1'b0};
7187: data_out = {8'd196, 8'd253, 1'b1, 1'b0};
7188: data_out = {8'd192, 8'd254, 1'b1, 1'b0};
7189: data_out = {8'd193, 8'd254, 1'b1, 1'b0};
7190: data_out = {8'd194, 8'd254, 1'b1, 1'b0};
7191: data_out = {8'd195, 8'd254, 1'b1, 1'b0};
7192: data_out = {8'd196, 8'd254, 1'b1, 1'b1};  //reset


            default: data_out = '0;
        endcase
    end

endmodule
