//////////////////////////////////////////////////////////////////////////////
/*
 Module name:   start_screen_rom
 Author:        kszdom, IG
 Description:   ROM memory for starting screen


  _   _ _    _  _____ _      ______          _____                        
 | \ | | |  | |/ ____| |    |  ____|   /\   |  __ \                       
 |  \| | |  | | |    | |    | |__     /  \  | |__) |                      
 | . ` | |  | | |    | |    |  __|   / /\ \ |  _  /                       
 | |\  | |__| | |____| |____| |____ / ____ \| | \ \                       
 |_| \_|\____/_\_____|______|______/_/_ __\_\_|__\_\  _____   ____  _   _ 
     /\   |  __ \|  \/  |   /\   / ____|  ____|  __ \|  __ \ / __ \| \ | |
    /  \  | |__) | \  / |  /  \ | |  __| |__  | |  | | |  | | |  | |  \| |
   / /\ \ |  _  /| |\/| | / /\ \| | |_ |  __| | |  | | |  | | |  | | . ` |
  / ____ \| | \ \| |  | |/ ____ \ |__| | |____| |__| | |__| | |__| | |\  |
 /_/___ \_\_|_ \_\_| _|_/_/__  \_\_____|______|_____/|_____/ \____/|_| \_|
 |_   _|/ ____| | \ | |  ____|   /\   |  __ \                             
   | | | (___   |  \| | |__     /  \  | |__) |                            
   | |  \___ \  | . ` |  __|   / /\ \ |  _  /                             
  _| |_ ____) | | |\  | |____ / ____ \| | \ \                             
 |_____|_____/  |_| \_|______/_/    \_\_|  \_\ 

 */
//////////////////////////////////////////////////////////////////////////////



module start_screen_rom #(
    parameter int ADDRESSWIDTH = 14,  // 4 bits => 16 entries
    parameter int DATAWIDTH = 18  // 8+8+1+1 = 18 bits
)(
    input logic [ADDRESSWIDTH-1:0] addr,
    output logic [DATAWIDTH-1:0] data_out
);


    always_comb begin
        unique case (addr)

            0: data_out = {8'd13, 8'd51, 1'b0, 1'b1};
            1: data_out = {8'd21, 8'd51, 1'b1, 1'b0};
            2: data_out = {8'd21, 8'd53, 1'b1, 1'b0};
            3: data_out = {8'd13, 8'd53, 1'b1, 1'b0};
            4: data_out = {8'd13, 8'd51, 1'b1, 1'b0};
            5: data_out = {8'd22, 8'd54, 1'b0, 1'b1};
            6: data_out = {8'd24, 8'd54, 1'b1, 1'b0};
            7: data_out = {8'd24, 8'd56, 1'b1, 1'b0};
            8: data_out = {8'd22, 8'd56, 1'b1, 1'b0};
            9: data_out = {8'd22, 8'd54, 1'b1, 1'b0};
            10: data_out = {8'd21, 8'd57, 1'b0, 1'b1};
            11: data_out = {8'd21, 8'd59, 1'b1, 1'b0};
            12: data_out = {8'd16, 8'd59, 1'b1, 1'b0};
            13: data_out = {8'd16, 8'd57, 1'b1, 1'b0};
            14: data_out = {8'd21, 8'd57, 1'b1, 1'b0};
            15: data_out = {8'd15, 8'd60, 1'b0, 1'b1};
            16: data_out = {8'd15, 8'd62, 1'b1, 1'b0};
            17: data_out = {8'd13, 8'd62, 1'b1, 1'b0};
            18: data_out = {8'd13, 8'd60, 1'b1, 1'b0};
            19: data_out = {8'd15, 8'd60, 1'b1, 1'b0};
            20: data_out = {8'd16, 8'd63, 1'b0, 1'b1};
            21: data_out = {8'd24, 8'd63, 1'b1, 1'b0};
            22: data_out = {8'd24, 8'd65, 1'b1, 1'b0};
            23: data_out = {8'd16, 8'd65, 1'b1, 1'b0};
            24: data_out = {8'd16, 8'd63, 1'b1, 1'b0};
            25: data_out = {8'd28, 8'd51, 1'b0, 1'b1};
            26: data_out = {8'd30, 8'd51, 1'b1, 1'b0};
            27: data_out = {8'd30, 8'd65, 1'b1, 1'b0};
            28: data_out = {8'd28, 8'd65, 1'b1, 1'b0};
            29: data_out = {8'd28, 8'd51, 1'b1, 1'b0};
            30: data_out = {8'd30, 8'd54, 1'b0, 1'b1};
            31: data_out = {8'd33, 8'd54, 1'b1, 1'b0};
            32: data_out = {8'd33, 8'd56, 1'b1, 1'b0};
            33: data_out = {8'd30, 8'd56, 1'b1, 1'b0};
            34: data_out = {8'd34, 8'd57, 1'b0, 1'b1};
            35: data_out = {8'd36, 8'd57, 1'b1, 1'b0};
            36: data_out = {8'd36, 8'd59, 1'b1, 1'b0};
            37: data_out = {8'd34, 8'd59, 1'b1, 1'b0};
            38: data_out = {8'd34, 8'd57, 1'b1, 1'b0};
            39: data_out = {8'd40, 8'd51, 1'b0, 1'b1};
            40: data_out = {8'd42, 8'd51, 1'b1, 1'b0};
            41: data_out = {8'd42, 8'd65, 1'b1, 1'b0};
            42: data_out = {8'd40, 8'd65, 1'b1, 1'b0};
            43: data_out = {8'd40, 8'd51, 1'b1, 1'b0};
            44: data_out = {8'd40, 8'd54, 1'b0, 1'b1};
            45: data_out = {8'd37, 8'd54, 1'b1, 1'b0};
            46: data_out = {8'd37, 8'd56, 1'b1, 1'b0};
            47: data_out = {8'd40, 8'd56, 1'b1, 1'b0};
            48: data_out = {8'd46, 8'd51, 1'b0, 1'b1};
            49: data_out = {8'd54, 8'd51, 1'b1, 1'b0};
            50: data_out = {8'd54, 8'd53, 1'b1, 1'b0};
            51: data_out = {8'd46, 8'd53, 1'b1, 1'b0};
            52: data_out = {8'd46, 8'd51, 1'b1, 1'b0};
            53: data_out = {8'd46, 8'd63, 1'b0, 1'b1};
            54: data_out = {8'd46, 8'd65, 1'b1, 1'b0};
            55: data_out = {8'd54, 8'd65, 1'b1, 1'b0};
            56: data_out = {8'd54, 8'd63, 1'b1, 1'b0};
            57: data_out = {8'd46, 8'd63, 1'b1, 1'b0};
            58: data_out = {8'd49, 8'd53, 1'b0, 1'b1};
            59: data_out = {8'd49, 8'd63, 1'b1, 1'b0};
            60: data_out = {8'd51, 8'd53, 1'b0, 1'b1};
            61: data_out = {8'd51, 8'd63, 1'b1, 1'b0};
            62: data_out = {8'd58, 8'd63, 1'b0, 1'b1};
            63: data_out = {8'd72, 8'd63, 1'b1, 1'b0};
            64: data_out = {8'd72, 8'd65, 1'b1, 1'b0};
            65: data_out = {8'd58, 8'd65, 1'b1, 1'b0};
            66: data_out = {8'd58, 8'd63, 1'b1, 1'b0};
            67: data_out = {8'd64, 8'd63, 1'b0, 1'b1};
            68: data_out = {8'd64, 8'd51, 1'b1, 1'b0};
            69: data_out = {8'd66, 8'd51, 1'b1, 1'b0};
            70: data_out = {8'd66, 8'd63, 1'b1, 1'b0};
            71: data_out = {8'd76, 8'd54, 1'b0, 1'b1};
            72: data_out = {8'd78, 8'd54, 1'b1, 1'b0};
            73: data_out = {8'd78, 8'd62, 1'b1, 1'b0};
            74: data_out = {8'd76, 8'd62, 1'b1, 1'b0};
            75: data_out = {8'd76, 8'd54, 1'b1, 1'b0};
            76: data_out = {8'd79, 8'd51, 1'b0, 1'b1};
            77: data_out = {8'd84, 8'd51, 1'b1, 1'b0};
            78: data_out = {8'd84, 8'd53, 1'b1, 1'b0};
            79: data_out = {8'd79, 8'd53, 1'b1, 1'b0};
            80: data_out = {8'd79, 8'd51, 1'b1, 1'b0};
            81: data_out = {8'd85, 8'd54, 1'b0, 1'b1};
            82: data_out = {8'd87, 8'd54, 1'b1, 1'b0};
            83: data_out = {8'd87, 8'd56, 1'b1, 1'b0};
            84: data_out = {8'd85, 8'd56, 1'b1, 1'b0};
            85: data_out = {8'd85, 8'd54, 1'b1, 1'b0};
            86: data_out = {8'd85, 8'd60, 1'b0, 1'b1};
            87: data_out = {8'd87, 8'd60, 1'b1, 1'b0};
            88: data_out = {8'd87, 8'd62, 1'b1, 1'b0};
            89: data_out = {8'd85, 8'd62, 1'b1, 1'b0};
            90: data_out = {8'd85, 8'd60, 1'b1, 1'b0};
            91: data_out = {8'd79, 8'd63, 1'b0, 1'b1};
            92: data_out = {8'd84, 8'd63, 1'b1, 1'b0};
            93: data_out = {8'd84, 8'd65, 1'b1, 1'b0};
            94: data_out = {8'd79, 8'd65, 1'b1, 1'b0};
            95: data_out = {8'd79, 8'd63, 1'b1, 1'b0};
            96: data_out = {8'd91, 8'd51, 1'b0, 1'b1};
            97: data_out = {8'd93, 8'd51, 1'b1, 1'b0};
            98: data_out = {8'd93, 8'd65, 1'b1, 1'b0};
            99: data_out = {8'd91, 8'd65, 1'b1, 1'b0};
            100: data_out = {8'd91, 8'd51, 1'b1, 1'b0};
            101: data_out = {8'd100, 8'd51, 1'b0, 1'b1};
            102: data_out = {8'd102, 8'd51, 1'b1, 1'b0};
            103: data_out = {8'd102, 8'd65, 1'b1, 1'b0};
            104: data_out = {8'd100, 8'd65, 1'b1, 1'b0};
            105: data_out = {8'd100, 8'd51, 1'b1, 1'b0};
            106: data_out = {8'd100, 8'd57, 1'b0, 1'b1};
            107: data_out = {8'd93, 8'd57, 1'b1, 1'b0};
            108: data_out = {8'd93, 8'd59, 1'b0, 1'b1};
            109: data_out = {8'd100, 8'd59, 1'b1, 1'b0};
            110: data_out = {8'd114, 8'd51, 1'b0, 1'b1};
            111: data_out = {8'd122, 8'd51, 1'b1, 1'b0};
            112: data_out = {8'd122, 8'd53, 1'b1, 1'b0};
            113: data_out = {8'd114, 8'd53, 1'b1, 1'b0};
            114: data_out = {8'd114, 8'd51, 1'b1, 1'b0};
            115: data_out = {8'd117, 8'd53, 1'b0, 1'b1};
            116: data_out = {8'd117, 8'd65, 1'b1, 1'b0};
            117: data_out = {8'd119, 8'd65, 1'b1, 1'b0};
            118: data_out = {8'd119, 8'd53, 1'b1, 1'b0};
            119: data_out = {8'd117, 8'd62, 1'b0, 1'b1};
            120: data_out = {8'd114, 8'd62, 1'b1, 1'b0};
            121: data_out = {8'd114, 8'd60, 1'b1, 1'b0};
            122: data_out = {8'd117, 8'd60, 1'b1, 1'b0};
            123: data_out = {8'd126, 8'd51, 1'b0, 1'b1};
            124: data_out = {8'd134, 8'd51, 1'b1, 1'b0};
            125: data_out = {8'd134, 8'd53, 1'b1, 1'b0};
            126: data_out = {8'd126, 8'd53, 1'b1, 1'b0};
            127: data_out = {8'd126, 8'd51, 1'b1, 1'b0};
            128: data_out = {8'd135, 8'd54, 1'b0, 1'b1};
            129: data_out = {8'd137, 8'd54, 1'b1, 1'b0};
            130: data_out = {8'd137, 8'd56, 1'b1, 1'b0};
            131: data_out = {8'd135, 8'd56, 1'b1, 1'b0};
            132: data_out = {8'd135, 8'd54, 1'b1, 1'b0};
            133: data_out = {8'd126, 8'd57, 1'b0, 1'b1};
            134: data_out = {8'd128, 8'd57, 1'b1, 1'b0};
            135: data_out = {8'd128, 8'd65, 1'b1, 1'b0};
            136: data_out = {8'd126, 8'd65, 1'b1, 1'b0};
            137: data_out = {8'd126, 8'd57, 1'b1, 1'b0};
            138: data_out = {8'd128, 8'd57, 1'b0, 1'b1};
            139: data_out = {8'd134, 8'd57, 1'b1, 1'b0};
            140: data_out = {8'd134, 8'd59, 1'b1, 1'b0};
            141: data_out = {8'd128, 8'd59, 1'b1, 1'b0};
            142: data_out = {8'd128, 8'd63, 1'b0, 1'b1};
            143: data_out = {8'd137, 8'd63, 1'b1, 1'b0};
            144: data_out = {8'd137, 8'd65, 1'b1, 1'b0};
            145: data_out = {8'd128, 8'd65, 1'b1, 1'b0};
            146: data_out = {8'd144, 8'd63, 1'b0, 1'b1};
            147: data_out = {8'd158, 8'd63, 1'b1, 1'b0};
            148: data_out = {8'd158, 8'd65, 1'b1, 1'b0};
            149: data_out = {8'd144, 8'd65, 1'b1, 1'b0};
            150: data_out = {8'd144, 8'd63, 1'b1, 1'b0};
            151: data_out = {8'd150, 8'd63, 1'b0, 1'b1};
            152: data_out = {8'd150, 8'd51, 1'b1, 1'b0};
            153: data_out = {8'd152, 8'd51, 1'b1, 1'b0};
            154: data_out = {8'd152, 8'd63, 1'b1, 1'b0};
            155: data_out = {8'd165, 8'd51, 1'b0, 1'b1};
            156: data_out = {8'd170, 8'd51, 1'b1, 1'b0};
            157: data_out = {8'd170, 8'd53, 1'b1, 1'b0};
            158: data_out = {8'd165, 8'd53, 1'b1, 1'b0};
            159: data_out = {8'd165, 8'd51, 1'b1, 1'b0};
            160: data_out = {8'd162, 8'd54, 1'b0, 1'b1};
            161: data_out = {8'd164, 8'd54, 1'b1, 1'b0};
            162: data_out = {8'd164, 8'd62, 1'b1, 1'b0};
            163: data_out = {8'd162, 8'd62, 1'b1, 1'b0};
            164: data_out = {8'd162, 8'd54, 1'b1, 1'b0};
            165: data_out = {8'd165, 8'd63, 1'b0, 1'b1};
            166: data_out = {8'd170, 8'd63, 1'b1, 1'b0};
            167: data_out = {8'd170, 8'd65, 1'b1, 1'b0};
            168: data_out = {8'd165, 8'd65, 1'b1, 1'b0};
            169: data_out = {8'd165, 8'd63, 1'b1, 1'b0};
            170: data_out = {8'd171, 8'd54, 1'b0, 1'b1};
            171: data_out = {8'd173, 8'd54, 1'b1, 1'b0};
            172: data_out = {8'd173, 8'd62, 1'b1, 1'b0};
            173: data_out = {8'd171, 8'd62, 1'b1, 1'b0};
            174: data_out = {8'd171, 8'd54, 1'b1, 1'b0};
            175: data_out = {8'd183, 8'd51, 1'b0, 1'b1};
            176: data_out = {8'd185, 8'd51, 1'b1, 1'b0};
            177: data_out = {8'd185, 8'd65, 1'b1, 1'b0};
            178: data_out = {8'd183, 8'd65, 1'b1, 1'b0};
            179: data_out = {8'd183, 8'd51, 1'b1, 1'b0};
            180: data_out = {8'd192, 8'd60, 1'b0, 1'b1};
            181: data_out = {8'd194, 8'd60, 1'b1, 1'b0};
            182: data_out = {8'd194, 8'd62, 1'b1, 1'b0};
            183: data_out = {8'd192, 8'd62, 1'b1, 1'b0};
            184: data_out = {8'd192, 8'd60, 1'b1, 1'b0};
            185: data_out = {8'd185, 8'd57, 1'b0, 1'b1};
            186: data_out = {8'd191, 8'd57, 1'b1, 1'b0};
            187: data_out = {8'd191, 8'd59, 1'b1, 1'b0};
            188: data_out = {8'd185, 8'd59, 1'b1, 1'b0};
            189: data_out = {8'd185, 8'd63, 1'b0, 1'b1};
            190: data_out = {8'd191, 8'd63, 1'b1, 1'b0};
            191: data_out = {8'd191, 8'd65, 1'b1, 1'b0};
            192: data_out = {8'd185, 8'd65, 1'b1, 1'b0};
            193: data_out = {8'd198, 8'd51, 1'b0, 1'b1};
            194: data_out = {8'd200, 8'd51, 1'b1, 1'b0};
            195: data_out = {8'd200, 8'd65, 1'b1, 1'b0};
            196: data_out = {8'd198, 8'd65, 1'b1, 1'b0};
            197: data_out = {8'd198, 8'd51, 1'b1, 1'b0};
            198: data_out = {8'd200, 8'd51, 1'b0, 1'b1};
            199: data_out = {8'd209, 8'd51, 1'b1, 1'b0};
            200: data_out = {8'd209, 8'd53, 1'b1, 1'b0};
            201: data_out = {8'd200, 8'd53, 1'b1, 1'b0};
            202: data_out = {8'd213, 8'd51, 1'b0, 1'b1};
            203: data_out = {8'd215, 8'd51, 1'b1, 1'b0};
            204: data_out = {8'd215, 8'd62, 1'b1, 1'b0};
            205: data_out = {8'd213, 8'd62, 1'b1, 1'b0};
            206: data_out = {8'd213, 8'd51, 1'b1, 1'b0};
            207: data_out = {8'd216, 8'd63, 1'b0, 1'b1};
            208: data_out = {8'd221, 8'd63, 1'b1, 1'b0};
            209: data_out = {8'd221, 8'd65, 1'b1, 1'b0};
            210: data_out = {8'd216, 8'd65, 1'b1, 1'b0};
            211: data_out = {8'd216, 8'd63, 1'b1, 1'b0};
            212: data_out = {8'd222, 8'd51, 1'b0, 1'b1};
            213: data_out = {8'd224, 8'd51, 1'b1, 1'b0};
            214: data_out = {8'd224, 8'd62, 1'b1, 1'b0};
            215: data_out = {8'd222, 8'd62, 1'b1, 1'b0};
            216: data_out = {8'd222, 8'd51, 1'b1, 1'b0};
            217: data_out = {8'd215, 8'd57, 1'b0, 1'b1};
            218: data_out = {8'd222, 8'd57, 1'b1, 1'b0};
            219: data_out = {8'd215, 8'd59, 1'b0, 1'b1};
            220: data_out = {8'd222, 8'd59, 1'b1, 1'b0};
            221: data_out = {8'd228, 8'd60, 1'b0, 1'b1};
            222: data_out = {8'd230, 8'd60, 1'b1, 1'b0};
            223: data_out = {8'd230, 8'd65, 1'b1, 1'b0};
            224: data_out = {8'd228, 8'd65, 1'b1, 1'b0};
            225: data_out = {8'd228, 8'd60, 1'b1, 1'b0};
            226: data_out = {8'd231, 8'd57, 1'b0, 1'b1};
            227: data_out = {8'd239, 8'd57, 1'b1, 1'b0};
            228: data_out = {8'd239, 8'd59, 1'b1, 1'b0};
            229: data_out = {8'd231, 8'd59, 1'b1, 1'b0};
            230: data_out = {8'd231, 8'd57, 1'b1, 1'b0};
            231: data_out = {8'd240, 8'd60, 1'b0, 1'b1};
            232: data_out = {8'd242, 8'd60, 1'b1, 1'b0};
            233: data_out = {8'd242, 8'd65, 1'b1, 1'b0};
            234: data_out = {8'd240, 8'd65, 1'b1, 1'b0};
            235: data_out = {8'd240, 8'd60, 1'b1, 1'b0};
            236: data_out = {8'd234, 8'd57, 1'b0, 1'b1};
            237: data_out = {8'd234, 8'd51, 1'b1, 1'b0};
            238: data_out = {8'd236, 8'd51, 1'b1, 1'b0};
            239: data_out = {8'd236, 8'd57, 1'b1, 1'b0};
            240: data_out = {8'd110, 8'd88, 1'b0, 1'b1};
            241: data_out = {8'd158, 8'd88, 1'b1, 1'b0};
            242: data_out = {8'd138, 8'd125, 1'b1, 1'b0};
            243: data_out = {8'd129, 8'd125, 1'b1, 1'b0};
            244: data_out = {8'd110, 8'd88, 1'b1, 1'b0};
            245: data_out = {8'd85, 8'd133, 1'b0, 1'b1};
            246: data_out = {8'd125, 8'd133, 1'b1, 1'b0};
            247: data_out = {8'd130, 8'd140, 1'b1, 1'b0};
            248: data_out = {8'd108, 8'd177, 1'b1, 1'b0};
            249: data_out = {8'd85, 8'd133, 1'b1, 1'b0};
            250: data_out = {8'd182, 8'd133, 1'b0, 1'b1};
            251: data_out = {8'd158, 8'd177, 1'b1, 1'b0};
            252: data_out = {8'd137, 8'd140, 1'b1, 1'b0};
            253: data_out = {8'd140, 8'd133, 1'b1, 1'b0};
            254: data_out = {8'd182, 8'd133, 1'b1, 1'b0};
            255: data_out = {8'd132, 8'd129, 1'b0, 1'b1};
            256: data_out = {8'd134, 8'd129, 1'b1, 1'b0};
            257: data_out = {8'd136, 8'd131, 1'b1, 1'b0};
            258: data_out = {8'd136, 8'd135, 1'b1, 1'b0};
            259: data_out = {8'd134, 8'd137, 1'b1, 1'b0};
            260: data_out = {8'd132, 8'd137, 1'b1, 1'b0};
            261: data_out = {8'd130, 8'd135, 1'b1, 1'b0};
            262: data_out = {8'd130, 8'd131, 1'b1, 1'b0};
            263: data_out = {8'd132, 8'd129, 1'b1, 1'b0};
            264: data_out = {8'd26, 8'd196, 1'b0, 1'b1};
            265: data_out = {8'd32, 8'd196, 1'b1, 1'b0};
            266: data_out = {8'd32, 8'd230, 1'b1, 1'b0};
            267: data_out = {8'd26, 8'd230, 1'b1, 1'b0};
            268: data_out = {8'd26, 8'd196, 1'b1, 1'b0};
            269: data_out = {8'd47, 8'd196, 1'b0, 1'b1};
            270: data_out = {8'd53, 8'd196, 1'b1, 1'b0};
            271: data_out = {8'd53, 8'd230, 1'b1, 1'b0};
            272: data_out = {8'd47, 8'd230, 1'b1, 1'b0};
            273: data_out = {8'd47, 8'd196, 1'b1, 1'b0};
            274: data_out = {8'd47, 8'd210, 1'b0, 1'b1};
            275: data_out = {8'd40, 8'd210, 1'b1, 1'b0};
            276: data_out = {8'd40, 8'd216, 1'b1, 1'b0};
            277: data_out = {8'd47, 8'd216, 1'b1, 1'b0};
            278: data_out = {8'd32, 8'd217, 1'b0, 1'b1};
            279: data_out = {8'd39, 8'd217, 1'b1, 1'b0};
            280: data_out = {8'd39, 8'd223, 1'b1, 1'b0};
            281: data_out = {8'd32, 8'd223, 1'b1, 1'b0};
            282: data_out = {8'd68, 8'd196, 1'b0, 1'b1};
            283: data_out = {8'd81, 8'd196, 1'b1, 1'b0};
            284: data_out = {8'd81, 8'd202, 1'b1, 1'b0};
            285: data_out = {8'd68, 8'd202, 1'b1, 1'b0};
            286: data_out = {8'd68, 8'd196, 1'b1, 1'b0};
            287: data_out = {8'd61, 8'd203, 1'b0, 1'b1};
            288: data_out = {8'd67, 8'd203, 1'b1, 1'b0};
            289: data_out = {8'd67, 8'd223, 1'b1, 1'b0};
            290: data_out = {8'd61, 8'd223, 1'b1, 1'b0};
            291: data_out = {8'd61, 8'd203, 1'b1, 1'b0};
            292: data_out = {8'd68, 8'd224, 1'b0, 1'b1};
            293: data_out = {8'd81, 8'd224, 1'b1, 1'b0};
            294: data_out = {8'd81, 8'd230, 1'b1, 1'b0};
            295: data_out = {8'd68, 8'd230, 1'b1, 1'b0};
            296: data_out = {8'd68, 8'd224, 1'b1, 1'b0};
            297: data_out = {8'd82, 8'd203, 1'b0, 1'b1};
            298: data_out = {8'd88, 8'd203, 1'b1, 1'b0};
            299: data_out = {8'd88, 8'd223, 1'b1, 1'b0};
            300: data_out = {8'd82, 8'd223, 1'b1, 1'b0};
            301: data_out = {8'd82, 8'd203, 1'b1, 1'b0};
            302: data_out = {8'd96, 8'd224, 1'b0, 1'b1};
            303: data_out = {8'd116, 8'd224, 1'b1, 1'b0};
            304: data_out = {8'd116, 8'd230, 1'b1, 1'b0};
            305: data_out = {8'd96, 8'd230, 1'b1, 1'b0};
            306: data_out = {8'd96, 8'd224, 1'b1, 1'b0};
            307: data_out = {8'd102, 8'd224, 1'b0, 1'b1};
            308: data_out = {8'd102, 8'd196, 1'b1, 1'b0};
            309: data_out = {8'd96, 8'd196, 1'b1, 1'b0};
            310: data_out = {8'd96, 8'd230, 1'b1, 1'b0};
            311: data_out = {8'd102, 8'd210, 1'b0, 1'b1};
            312: data_out = {8'd116, 8'd210, 1'b1, 1'b0};
            313: data_out = {8'd116, 8'd216, 1'b1, 1'b0};
            314: data_out = {8'd102, 8'd216, 1'b1, 1'b0};
            315: data_out = {8'd117, 8'd217, 1'b0, 1'b1};
            316: data_out = {8'd123, 8'd217, 1'b1, 1'b0};
            317: data_out = {8'd123, 8'd223, 1'b1, 1'b0};
            318: data_out = {8'd117, 8'd223, 1'b1, 1'b0};
            319: data_out = {8'd117, 8'd217, 1'b1, 1'b0};
            320: data_out = {8'd117, 8'd196, 1'b0, 1'b1};
            321: data_out = {8'd123, 8'd196, 1'b1, 1'b0};
            322: data_out = {8'd123, 8'd202, 1'b1, 1'b0};
            323: data_out = {8'd117, 8'd202, 1'b1, 1'b0};
            324: data_out = {8'd117, 8'd196, 1'b1, 1'b0};
            325: data_out = {8'd110, 8'd210, 1'b0, 1'b1};
            326: data_out = {8'd110, 8'd203, 1'b1, 1'b0};
            327: data_out = {8'd116, 8'd203, 1'b1, 1'b0};
            328: data_out = {8'd116, 8'd210, 1'b1, 1'b0};
            329: data_out = {8'd131, 8'd196, 1'b0, 1'b1};
            330: data_out = {8'd137, 8'd196, 1'b1, 1'b0};
            331: data_out = {8'd137, 8'd223, 1'b1, 1'b0};
            332: data_out = {8'd131, 8'd223, 1'b1, 1'b0};
            333: data_out = {8'd131, 8'd196, 1'b1, 1'b0};
            334: data_out = {8'd152, 8'd196, 1'b0, 1'b1};
            335: data_out = {8'd158, 8'd196, 1'b1, 1'b0};
            336: data_out = {8'd158, 8'd223, 1'b1, 1'b0};
            337: data_out = {8'd152, 8'd223, 1'b1, 1'b0};
            338: data_out = {8'd152, 8'd196, 1'b1, 1'b0};
            339: data_out = {8'd138, 8'd224, 1'b0, 1'b1};
            340: data_out = {8'd151, 8'd224, 1'b1, 1'b0};
            341: data_out = {8'd151, 8'd230, 1'b1, 1'b0};
            342: data_out = {8'd138, 8'd230, 1'b1, 1'b0};
            343: data_out = {8'd138, 8'd224, 1'b1, 1'b0};
            344: data_out = {8'd137, 8'd210, 1'b0, 1'b1};
            345: data_out = {8'd152, 8'd210, 1'b1, 1'b0};
            346: data_out = {8'd137, 8'd216, 1'b0, 1'b1};
            347: data_out = {8'd152, 8'd216, 1'b1, 1'b0};
            348: data_out = {8'd166, 8'd196, 1'b0, 1'b1};
            349: data_out = {8'd186, 8'd196, 1'b1, 1'b0};
            350: data_out = {8'd186, 8'd202, 1'b1, 1'b0};
            351: data_out = {8'd166, 8'd202, 1'b1, 1'b0};
            352: data_out = {8'd166, 8'd196, 1'b1, 1'b0};
            353: data_out = {8'd166, 8'd224, 1'b0, 1'b1};
            354: data_out = {8'd186, 8'd224, 1'b1, 1'b0};
            355: data_out = {8'd186, 8'd230, 1'b1, 1'b0};
            356: data_out = {8'd166, 8'd230, 1'b1, 1'b0};
            357: data_out = {8'd166, 8'd224, 1'b1, 1'b0};
            358: data_out = {8'd187, 8'd203, 1'b0, 1'b1};
            359: data_out = {8'd193, 8'd203, 1'b1, 1'b0};
            360: data_out = {8'd193, 8'd223, 1'b1, 1'b0};
            361: data_out = {8'd187, 8'd223, 1'b1, 1'b0};
            362: data_out = {8'd187, 8'd203, 1'b1, 1'b0};
            363: data_out = {8'd166, 8'd202, 1'b0, 1'b1};
            364: data_out = {8'd166, 8'd224, 1'b1, 1'b0};
            365: data_out = {8'd172, 8'd202, 1'b0, 1'b1};
            366: data_out = {8'd172, 8'd224, 1'b1, 1'b0};
            367: data_out = {8'd198, 8'd210, 1'b0, 1'b1};
            368: data_out = {8'd210, 8'd210, 1'b1, 1'b0};
            369: data_out = {8'd210, 8'd216, 1'b1, 1'b0};
            370: data_out = {8'd198, 8'd216, 1'b1, 1'b0};
            371: data_out = {8'd198, 8'd210, 1'b1, 1'b0};
            372: data_out = {8'd215, 8'd196, 1'b0, 1'b1};
            373: data_out = {8'd221, 8'd196, 1'b1, 1'b0};
            374: data_out = {8'd221, 8'd223, 1'b1, 1'b0};
            375: data_out = {8'd215, 8'd223, 1'b1, 1'b0};
            376: data_out = {8'd215, 8'd196, 1'b1, 1'b0};
            377: data_out = {8'd236, 8'd196, 1'b0, 1'b1};
            378: data_out = {8'd242, 8'd196, 1'b1, 1'b0};
            379: data_out = {8'd242, 8'd223, 1'b1, 1'b0};
            380: data_out = {8'd236, 8'd223, 1'b1, 1'b0};
            381: data_out = {8'd236, 8'd196, 1'b1, 1'b0};
            382: data_out = {8'd222, 8'd224, 1'b0, 1'b1};
            383: data_out = {8'd235, 8'd224, 1'b1, 1'b0};
            384: data_out = {8'd235, 8'd230, 1'b1, 1'b0};
            385: data_out = {8'd222, 8'd230, 1'b1, 1'b0};
            386: data_out = {8'd222, 8'd224, 1'b1, 1'b0};
            387: data_out = {8'd221, 8'd210, 1'b0, 1'b1};
            388: data_out = {8'd236, 8'd210, 1'b1, 1'b0};
            389: data_out = {8'd221, 8'd216, 1'b0, 1'b1};
            390: data_out = {8'd236, 8'd216, 1'b1, 1'b0};
            391: data_out = {8'd236, 8'd216, 1'b1, 1'b1};

            default: data_out = {8'd0, 8'd0, 1'b1, 1'b1};
        endcase
    end

endmodule
