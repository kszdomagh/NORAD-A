//////////////////////////////////////////////////////////////////////////////
/*
 Module name:   ending_screen_rom
 Author:        kszdom
 Description:   ROM memory for ending screen


  _   _ _    _  _____ _      ______          _____                        
 | \ | | |  | |/ ____| |    |  ____|   /\   |  __ \                       
 |  \| | |  | | |    | |    | |__     /  \  | |__) |                      
 | . ` | |  | | |    | |    |  __|   / /\ \ |  _  /                       
 | |\  | |__| | |____| |____| |____ / ____ \| | \ \                       
 |_| \_|\____/_\_____|______|______/_/_ __\_\_|__\_\  _____   ____  _   _ 
     /\   |  __ \|  \/  |   /\   / ____|  ____|  __ \|  __ \ / __ \| \ | |
    /  \  | |__) | \  / |  /  \ | |  __| |__  | |  | | |  | | |  | |  \| |
   / /\ \ |  _  /| |\/| | / /\ \| | |_ |  __| | |  | | |  | | |  | | . ` |
  / ____ \| | \ \| |  | |/ ____ \ |__| | |____| |__| | |__| | |__| | |\  |
 /_/___ \_\_|_ \_\_| _|_/_/__  \_\_____|______|_____/|_____/ \____/|_| \_|
 |_   _|/ ____| | \ | |  ____|   /\   |  __ \                             
   | | | (___   |  \| | |__     /  \  | |__) |                            
   | |  \___ \  | . ` |  __|   / /\ \ |  _  /                             
  _| |_ ____) | | |\  | |____ / ____ \| | \ \                             
 |_____|_____/  |_| \_|______/_/    \_\_|  \_\ 

 */
//////////////////////////////////////////////////////////////////////////////



module end_screen_rom #(
    parameter int ADDRESSWIDTH = 4,  // 4 bits => 16 entries
    parameter int DATAWIDTH = 18  // 8+8+1+1 = 18 bits
)(
    input logic [ADDRESSWIDTH-1:0] addr,
    output logic [DATAWIDTH-1:0] data_out
);

    always_comb begin
        unique case (addr)
            //                  x       y       line    pos

0: data_out = {8'd37, 8'd15, 1'b1, 1'b0};
1: data_out = {8'd38, 8'd15, 1'b1, 1'b0};
2: data_out = {8'd39, 8'd15, 1'b1, 1'b0};
3: data_out = {8'd40, 8'd15, 1'b1, 1'b0};
4: data_out = {8'd41, 8'd15, 1'b1, 1'b0};
5: data_out = {8'd42, 8'd15, 1'b1, 1'b0};
6: data_out = {8'd43, 8'd15, 1'b1, 1'b0};
7: data_out = {8'd44, 8'd15, 1'b1, 1'b0};
8: data_out = {8'd45, 8'd15, 1'b1, 1'b0};
9: data_out = {8'd46, 8'd15, 1'b1, 1'b0};
10: data_out = {8'd49, 8'd15, 1'b1, 1'b0};
11: data_out = {8'd50, 8'd15, 1'b1, 1'b0};
12: data_out = {8'd51, 8'd15, 1'b1, 1'b0};
13: data_out = {8'd52, 8'd15, 1'b1, 1'b0};
14: data_out = {8'd53, 8'd15, 1'b1, 1'b0};
15: data_out = {8'd54, 8'd15, 1'b1, 1'b0};
16: data_out = {8'd55, 8'd15, 1'b1, 1'b0};
17: data_out = {8'd56, 8'd15, 1'b1, 1'b0};
18: data_out = {8'd57, 8'd15, 1'b1, 1'b0};
19: data_out = {8'd58, 8'd15, 1'b1, 1'b0};
20: data_out = {8'd59, 8'd15, 1'b1, 1'b0};
21: data_out = {8'd60, 8'd15, 1'b1, 1'b0};
22: data_out = {8'd61, 8'd15, 1'b1, 1'b0};
23: data_out = {8'd62, 8'd15, 1'b1, 1'b0};
24: data_out = {8'd63, 8'd15, 1'b1, 1'b0};
25: data_out = {8'd64, 8'd15, 1'b1, 1'b0};
26: data_out = {8'd65, 8'd15, 1'b1, 1'b0};
27: data_out = {8'd66, 8'd15, 1'b1, 1'b0};
28: data_out = {8'd86, 8'd15, 1'b1, 1'b0};
29: data_out = {8'd87, 8'd15, 1'b1, 1'b0};
30: data_out = {8'd88, 8'd15, 1'b1, 1'b0};
31: data_out = {8'd89, 8'd15, 1'b1, 1'b0};
32: data_out = {8'd90, 8'd15, 1'b1, 1'b0};
33: data_out = {8'd91, 8'd15, 1'b1, 1'b0};
34: data_out = {8'd92, 8'd15, 1'b1, 1'b0};
35: data_out = {8'd93, 8'd15, 1'b1, 1'b0};
36: data_out = {8'd94, 8'd15, 1'b1, 1'b0};
37: data_out = {8'd95, 8'd15, 1'b1, 1'b0};
38: data_out = {8'd96, 8'd15, 1'b1, 1'b0};
39: data_out = {8'd97, 8'd15, 1'b1, 1'b0};
40: data_out = {8'd98, 8'd15, 1'b1, 1'b0};
41: data_out = {8'd99, 8'd15, 1'b1, 1'b0};
42: data_out = {8'd100, 8'd15, 1'b1, 1'b0};
43: data_out = {8'd101, 8'd15, 1'b1, 1'b0};
44: data_out = {8'd102, 8'd15, 1'b1, 1'b0};
45: data_out = {8'd103, 8'd15, 1'b1, 1'b0};
46: data_out = {8'd104, 8'd15, 1'b1, 1'b0};
47: data_out = {8'd105, 8'd15, 1'b1, 1'b0};
48: data_out = {8'd106, 8'd15, 1'b1, 1'b0};
49: data_out = {8'd107, 8'd15, 1'b1, 1'b0};
50: data_out = {8'd108, 8'd15, 1'b1, 1'b0};
51: data_out = {8'd109, 8'd15, 1'b1, 1'b0};
52: data_out = {8'd110, 8'd15, 1'b1, 1'b0};
53: data_out = {8'd111, 8'd15, 1'b1, 1'b0};
54: data_out = {8'd112, 8'd15, 1'b1, 1'b0};
55: data_out = {8'd113, 8'd15, 1'b1, 1'b0};
56: data_out = {8'd114, 8'd15, 1'b1, 1'b0};
57: data_out = {8'd115, 8'd15, 1'b1, 1'b0};
58: data_out = {8'd147, 8'd15, 1'b1, 1'b0};
59: data_out = {8'd148, 8'd15, 1'b1, 1'b0};
60: data_out = {8'd149, 8'd15, 1'b1, 1'b0};
61: data_out = {8'd150, 8'd15, 1'b1, 1'b0};
62: data_out = {8'd151, 8'd15, 1'b1, 1'b0};
63: data_out = {8'd152, 8'd15, 1'b1, 1'b0};
64: data_out = {8'd153, 8'd15, 1'b1, 1'b0};
65: data_out = {8'd154, 8'd15, 1'b1, 1'b0};
66: data_out = {8'd155, 8'd15, 1'b1, 1'b0};
67: data_out = {8'd156, 8'd15, 1'b1, 1'b0};
68: data_out = {8'd192, 8'd15, 1'b1, 1'b0};
69: data_out = {8'd193, 8'd15, 1'b1, 1'b0};
70: data_out = {8'd194, 8'd15, 1'b1, 1'b0};
71: data_out = {8'd195, 8'd15, 1'b1, 1'b0};
72: data_out = {8'd196, 8'd15, 1'b1, 1'b0};
73: data_out = {8'd197, 8'd15, 1'b1, 1'b0};
74: data_out = {8'd198, 8'd15, 1'b1, 1'b0};
75: data_out = {8'd199, 8'd15, 1'b1, 1'b0};
76: data_out = {8'd200, 8'd15, 1'b1, 1'b0};
77: data_out = {8'd201, 8'd15, 1'b1, 1'b0};
78: data_out = {8'd202, 8'd15, 1'b1, 1'b0};
79: data_out = {8'd203, 8'd15, 1'b1, 1'b0};
80: data_out = {8'd204, 8'd15, 1'b1, 1'b0};
81: data_out = {8'd205, 8'd15, 1'b1, 1'b0};
82: data_out = {8'd37, 8'd16, 1'b1, 1'b0};
83: data_out = {8'd46, 8'd16, 1'b1, 1'b0};
84: data_out = {8'd49, 8'd16, 1'b1, 1'b0};
85: data_out = {8'd66, 8'd16, 1'b1, 1'b0};
86: data_out = {8'd86, 8'd16, 1'b1, 1'b0};
87: data_out = {8'd115, 8'd16, 1'b1, 1'b0};
88: data_out = {8'd147, 8'd16, 1'b1, 1'b0};
89: data_out = {8'd156, 8'd16, 1'b1, 1'b0};
90: data_out = {8'd192, 8'd16, 1'b1, 1'b0};
91: data_out = {8'd205, 8'd16, 1'b1, 1'b0};
92: data_out = {8'd37, 8'd17, 1'b1, 1'b0};
93: data_out = {8'd46, 8'd17, 1'b1, 1'b0};
94: data_out = {8'd49, 8'd17, 1'b1, 1'b0};
95: data_out = {8'd66, 8'd17, 1'b1, 1'b0};
96: data_out = {8'd86, 8'd17, 1'b1, 1'b0};
97: data_out = {8'd115, 8'd17, 1'b1, 1'b0};
98: data_out = {8'd147, 8'd17, 1'b1, 1'b0};
99: data_out = {8'd156, 8'd17, 1'b1, 1'b0};
100: data_out = {8'd192, 8'd17, 1'b1, 1'b0};
101: data_out = {8'd205, 8'd17, 1'b1, 1'b0};
102: data_out = {8'd37, 8'd18, 1'b1, 1'b0};
103: data_out = {8'd46, 8'd18, 1'b1, 1'b0};
104: data_out = {8'd49, 8'd18, 1'b1, 1'b0};
105: data_out = {8'd66, 8'd18, 1'b1, 1'b0};
106: data_out = {8'd86, 8'd18, 1'b1, 1'b0};
107: data_out = {8'd115, 8'd18, 1'b1, 1'b0};
108: data_out = {8'd147, 8'd18, 1'b1, 1'b0};
109: data_out = {8'd156, 8'd18, 1'b1, 1'b0};
110: data_out = {8'd192, 8'd18, 1'b1, 1'b0};
111: data_out = {8'd205, 8'd18, 1'b1, 1'b0};
112: data_out = {8'd37, 8'd19, 1'b1, 1'b0};
113: data_out = {8'd46, 8'd19, 1'b1, 1'b0};
114: data_out = {8'd49, 8'd19, 1'b1, 1'b0};
115: data_out = {8'd50, 8'd19, 1'b1, 1'b0};
116: data_out = {8'd51, 8'd19, 1'b1, 1'b0};
117: data_out = {8'd52, 8'd19, 1'b1, 1'b0};
118: data_out = {8'd53, 8'd19, 1'b1, 1'b0};
119: data_out = {8'd62, 8'd19, 1'b1, 1'b0};
120: data_out = {8'd63, 8'd19, 1'b1, 1'b0};
121: data_out = {8'd64, 8'd19, 1'b1, 1'b0};
122: data_out = {8'd65, 8'd19, 1'b1, 1'b0};
123: data_out = {8'd66, 8'd19, 1'b1, 1'b0};
124: data_out = {8'd86, 8'd19, 1'b1, 1'b0};
125: data_out = {8'd91, 8'd19, 1'b1, 1'b0};
126: data_out = {8'd92, 8'd19, 1'b1, 1'b0};
127: data_out = {8'd93, 8'd19, 1'b1, 1'b0};
128: data_out = {8'd94, 8'd19, 1'b1, 1'b0};
129: data_out = {8'd95, 8'd19, 1'b1, 1'b0};
130: data_out = {8'd96, 8'd19, 1'b1, 1'b0};
131: data_out = {8'd97, 8'd19, 1'b1, 1'b0};
132: data_out = {8'd98, 8'd19, 1'b1, 1'b0};
133: data_out = {8'd99, 8'd19, 1'b1, 1'b0};
134: data_out = {8'd100, 8'd19, 1'b1, 1'b0};
135: data_out = {8'd101, 8'd19, 1'b1, 1'b0};
136: data_out = {8'd102, 8'd19, 1'b1, 1'b0};
137: data_out = {8'd111, 8'd19, 1'b1, 1'b0};
138: data_out = {8'd112, 8'd19, 1'b1, 1'b0};
139: data_out = {8'd113, 8'd19, 1'b1, 1'b0};
140: data_out = {8'd114, 8'd19, 1'b1, 1'b0};
141: data_out = {8'd115, 8'd19, 1'b1, 1'b0};
142: data_out = {8'd143, 8'd19, 1'b1, 1'b0};
143: data_out = {8'd144, 8'd19, 1'b1, 1'b0};
144: data_out = {8'd145, 8'd19, 1'b1, 1'b0};
145: data_out = {8'd146, 8'd19, 1'b1, 1'b0};
146: data_out = {8'd147, 8'd19, 1'b1, 1'b0};
147: data_out = {8'd156, 8'd19, 1'b1, 1'b0};
148: data_out = {8'd157, 8'd19, 1'b1, 1'b0};
149: data_out = {8'd158, 8'd19, 1'b1, 1'b0};
150: data_out = {8'd159, 8'd19, 1'b1, 1'b0};
151: data_out = {8'd160, 8'd19, 1'b1, 1'b0};
152: data_out = {8'd188, 8'd19, 1'b1, 1'b0};
153: data_out = {8'd189, 8'd19, 1'b1, 1'b0};
154: data_out = {8'd190, 8'd19, 1'b1, 1'b0};
155: data_out = {8'd191, 8'd19, 1'b1, 1'b0};
156: data_out = {8'd192, 8'd19, 1'b1, 1'b0};
157: data_out = {8'd197, 8'd19, 1'b1, 1'b0};
158: data_out = {8'd198, 8'd19, 1'b1, 1'b0};
159: data_out = {8'd199, 8'd19, 1'b1, 1'b0};
160: data_out = {8'd200, 8'd19, 1'b1, 1'b0};
161: data_out = {8'd205, 8'd19, 1'b1, 1'b0};
162: data_out = {8'd206, 8'd19, 1'b1, 1'b0};
163: data_out = {8'd207, 8'd19, 1'b1, 1'b0};
164: data_out = {8'd208, 8'd19, 1'b1, 1'b0};
165: data_out = {8'd209, 8'd19, 1'b1, 1'b0};
166: data_out = {8'd37, 8'd20, 1'b1, 1'b0};
167: data_out = {8'd46, 8'd20, 1'b1, 1'b0};
168: data_out = {8'd53, 8'd20, 1'b1, 1'b0};
169: data_out = {8'd62, 8'd20, 1'b1, 1'b0};
170: data_out = {8'd86, 8'd20, 1'b1, 1'b0};
171: data_out = {8'd91, 8'd20, 1'b1, 1'b0};
172: data_out = {8'd102, 8'd20, 1'b1, 1'b0};
173: data_out = {8'd111, 8'd20, 1'b1, 1'b0};
174: data_out = {8'd143, 8'd20, 1'b1, 1'b0};
175: data_out = {8'd160, 8'd20, 1'b1, 1'b0};
176: data_out = {8'd188, 8'd20, 1'b1, 1'b0};
177: data_out = {8'd197, 8'd20, 1'b1, 1'b0};
178: data_out = {8'd200, 8'd20, 1'b1, 1'b0};
179: data_out = {8'd209, 8'd20, 1'b1, 1'b0};
180: data_out = {8'd37, 8'd21, 1'b1, 1'b0};
181: data_out = {8'd46, 8'd21, 1'b1, 1'b0};
182: data_out = {8'd53, 8'd21, 1'b1, 1'b0};
183: data_out = {8'd62, 8'd21, 1'b1, 1'b0};
184: data_out = {8'd86, 8'd21, 1'b1, 1'b0};
185: data_out = {8'd91, 8'd21, 1'b1, 1'b0};
186: data_out = {8'd102, 8'd21, 1'b1, 1'b0};
187: data_out = {8'd111, 8'd21, 1'b1, 1'b0};
188: data_out = {8'd143, 8'd21, 1'b1, 1'b0};
189: data_out = {8'd160, 8'd21, 1'b1, 1'b0};
190: data_out = {8'd188, 8'd21, 1'b1, 1'b0};
191: data_out = {8'd197, 8'd21, 1'b1, 1'b0};
192: data_out = {8'd200, 8'd21, 1'b1, 1'b0};
193: data_out = {8'd209, 8'd21, 1'b1, 1'b0};
194: data_out = {8'd37, 8'd22, 1'b1, 1'b0};
195: data_out = {8'd46, 8'd22, 1'b1, 1'b0};
196: data_out = {8'd53, 8'd22, 1'b1, 1'b0};
197: data_out = {8'd62, 8'd22, 1'b1, 1'b0};
198: data_out = {8'd86, 8'd22, 1'b1, 1'b0};
199: data_out = {8'd91, 8'd22, 1'b1, 1'b0};
200: data_out = {8'd102, 8'd22, 1'b1, 1'b0};
201: data_out = {8'd111, 8'd22, 1'b1, 1'b0};
202: data_out = {8'd143, 8'd22, 1'b1, 1'b0};
203: data_out = {8'd160, 8'd22, 1'b1, 1'b0};
204: data_out = {8'd188, 8'd22, 1'b1, 1'b0};
205: data_out = {8'd197, 8'd22, 1'b1, 1'b0};
206: data_out = {8'd200, 8'd22, 1'b1, 1'b0};
207: data_out = {8'd209, 8'd22, 1'b1, 1'b0};
208: data_out = {8'd37, 8'd23, 1'b1, 1'b0};
209: data_out = {8'd46, 8'd23, 1'b1, 1'b0};
210: data_out = {8'd53, 8'd23, 1'b1, 1'b0};
211: data_out = {8'd62, 8'd23, 1'b1, 1'b0};
212: data_out = {8'd86, 8'd23, 1'b1, 1'b0};
213: data_out = {8'd87, 8'd23, 1'b1, 1'b0};
214: data_out = {8'd88, 8'd23, 1'b1, 1'b0};
215: data_out = {8'd89, 8'd23, 1'b1, 1'b0};
216: data_out = {8'd90, 8'd23, 1'b1, 1'b0};
217: data_out = {8'd91, 8'd23, 1'b1, 1'b0};
218: data_out = {8'd102, 8'd23, 1'b1, 1'b0};
219: data_out = {8'd111, 8'd23, 1'b1, 1'b0};
220: data_out = {8'd139, 8'd23, 1'b1, 1'b0};
221: data_out = {8'd140, 8'd23, 1'b1, 1'b0};
222: data_out = {8'd141, 8'd23, 1'b1, 1'b0};
223: data_out = {8'd142, 8'd23, 1'b1, 1'b0};
224: data_out = {8'd143, 8'd23, 1'b1, 1'b0};
225: data_out = {8'd148, 8'd23, 1'b1, 1'b0};
226: data_out = {8'd149, 8'd23, 1'b1, 1'b0};
227: data_out = {8'd150, 8'd23, 1'b1, 1'b0};
228: data_out = {8'd151, 8'd23, 1'b1, 1'b0};
229: data_out = {8'd152, 8'd23, 1'b1, 1'b0};
230: data_out = {8'd153, 8'd23, 1'b1, 1'b0};
231: data_out = {8'd154, 8'd23, 1'b1, 1'b0};
232: data_out = {8'd155, 8'd23, 1'b1, 1'b0};
233: data_out = {8'd160, 8'd23, 1'b1, 1'b0};
234: data_out = {8'd161, 8'd23, 1'b1, 1'b0};
235: data_out = {8'd162, 8'd23, 1'b1, 1'b0};
236: data_out = {8'd163, 8'd23, 1'b1, 1'b0};
237: data_out = {8'd164, 8'd23, 1'b1, 1'b0};
238: data_out = {8'd184, 8'd23, 1'b1, 1'b0};
239: data_out = {8'd185, 8'd23, 1'b1, 1'b0};
240: data_out = {8'd186, 8'd23, 1'b1, 1'b0};
241: data_out = {8'd187, 8'd23, 1'b1, 1'b0};
242: data_out = {8'd188, 8'd23, 1'b1, 1'b0};
243: data_out = {8'd193, 8'd23, 1'b1, 1'b0};
244: data_out = {8'd194, 8'd23, 1'b1, 1'b0};
245: data_out = {8'd195, 8'd23, 1'b1, 1'b0};
246: data_out = {8'd196, 8'd23, 1'b1, 1'b0};
247: data_out = {8'd197, 8'd23, 1'b1, 1'b0};
248: data_out = {8'd200, 8'd23, 1'b1, 1'b0};
249: data_out = {8'd201, 8'd23, 1'b1, 1'b0};
250: data_out = {8'd202, 8'd23, 1'b1, 1'b0};
251: data_out = {8'd203, 8'd23, 1'b1, 1'b0};
252: data_out = {8'd204, 8'd23, 1'b1, 1'b0};
253: data_out = {8'd209, 8'd23, 1'b1, 1'b0};
254: data_out = {8'd210, 8'd23, 1'b1, 1'b0};
255: data_out = {8'd211, 8'd23, 1'b1, 1'b0};
256: data_out = {8'd212, 8'd23, 1'b1, 1'b0};
257: data_out = {8'd213, 8'd23, 1'b1, 1'b0};
258: data_out = {8'd37, 8'd24, 1'b1, 1'b0};
259: data_out = {8'd46, 8'd24, 1'b1, 1'b0};
260: data_out = {8'd53, 8'd24, 1'b1, 1'b0};
261: data_out = {8'd62, 8'd24, 1'b1, 1'b0};
262: data_out = {8'd102, 8'd24, 1'b1, 1'b0};
263: data_out = {8'd111, 8'd24, 1'b1, 1'b0};
264: data_out = {8'd139, 8'd24, 1'b1, 1'b0};
265: data_out = {8'd148, 8'd24, 1'b1, 1'b0};
266: data_out = {8'd155, 8'd24, 1'b1, 1'b0};
267: data_out = {8'd164, 8'd24, 1'b1, 1'b0};
268: data_out = {8'd184, 8'd24, 1'b1, 1'b0};
269: data_out = {8'd193, 8'd24, 1'b1, 1'b0};
270: data_out = {8'd204, 8'd24, 1'b1, 1'b0};
271: data_out = {8'd213, 8'd24, 1'b1, 1'b0};
272: data_out = {8'd37, 8'd25, 1'b1, 1'b0};
273: data_out = {8'd46, 8'd25, 1'b1, 1'b0};
274: data_out = {8'd53, 8'd25, 1'b1, 1'b0};
275: data_out = {8'd62, 8'd25, 1'b1, 1'b0};
276: data_out = {8'd102, 8'd25, 1'b1, 1'b0};
277: data_out = {8'd111, 8'd25, 1'b1, 1'b0};
278: data_out = {8'd139, 8'd25, 1'b1, 1'b0};
279: data_out = {8'd148, 8'd25, 1'b1, 1'b0};
280: data_out = {8'd155, 8'd25, 1'b1, 1'b0};
281: data_out = {8'd164, 8'd25, 1'b1, 1'b0};
282: data_out = {8'd184, 8'd25, 1'b1, 1'b0};
283: data_out = {8'd193, 8'd25, 1'b1, 1'b0};
284: data_out = {8'd204, 8'd25, 1'b1, 1'b0};
285: data_out = {8'd213, 8'd25, 1'b1, 1'b0};
286: data_out = {8'd37, 8'd26, 1'b1, 1'b0};
287: data_out = {8'd46, 8'd26, 1'b1, 1'b0};
288: data_out = {8'd53, 8'd26, 1'b1, 1'b0};
289: data_out = {8'd62, 8'd26, 1'b1, 1'b0};
290: data_out = {8'd102, 8'd26, 1'b1, 1'b0};
291: data_out = {8'd111, 8'd26, 1'b1, 1'b0};
292: data_out = {8'd139, 8'd26, 1'b1, 1'b0};
293: data_out = {8'd148, 8'd26, 1'b1, 1'b0};
294: data_out = {8'd155, 8'd26, 1'b1, 1'b0};
295: data_out = {8'd164, 8'd26, 1'b1, 1'b0};
296: data_out = {8'd184, 8'd26, 1'b1, 1'b0};
297: data_out = {8'd193, 8'd26, 1'b1, 1'b0};
298: data_out = {8'd204, 8'd26, 1'b1, 1'b0};
299: data_out = {8'd213, 8'd26, 1'b1, 1'b0};
300: data_out = {8'd37, 8'd27, 1'b1, 1'b0};
301: data_out = {8'd38, 8'd27, 1'b1, 1'b0};
302: data_out = {8'd39, 8'd27, 1'b1, 1'b0};
303: data_out = {8'd40, 8'd27, 1'b1, 1'b0};
304: data_out = {8'd41, 8'd27, 1'b1, 1'b0};
305: data_out = {8'd46, 8'd27, 1'b1, 1'b0};
306: data_out = {8'd47, 8'd27, 1'b1, 1'b0};
307: data_out = {8'd48, 8'd27, 1'b1, 1'b0};
308: data_out = {8'd49, 8'd27, 1'b1, 1'b0};
309: data_out = {8'd50, 8'd27, 1'b1, 1'b0};
310: data_out = {8'd53, 8'd27, 1'b1, 1'b0};
311: data_out = {8'd62, 8'd27, 1'b1, 1'b0};
312: data_out = {8'd90, 8'd27, 1'b1, 1'b0};
313: data_out = {8'd91, 8'd27, 1'b1, 1'b0};
314: data_out = {8'd92, 8'd27, 1'b1, 1'b0};
315: data_out = {8'd93, 8'd27, 1'b1, 1'b0};
316: data_out = {8'd94, 8'd27, 1'b1, 1'b0};
317: data_out = {8'd95, 8'd27, 1'b1, 1'b0};
318: data_out = {8'd102, 8'd27, 1'b1, 1'b0};
319: data_out = {8'd111, 8'd27, 1'b1, 1'b0};
320: data_out = {8'd139, 8'd27, 1'b1, 1'b0};
321: data_out = {8'd148, 8'd27, 1'b1, 1'b0};
322: data_out = {8'd155, 8'd27, 1'b1, 1'b0};
323: data_out = {8'd164, 8'd27, 1'b1, 1'b0};
324: data_out = {8'd184, 8'd27, 1'b1, 1'b0};
325: data_out = {8'd193, 8'd27, 1'b1, 1'b0};
326: data_out = {8'd204, 8'd27, 1'b1, 1'b0};
327: data_out = {8'd213, 8'd27, 1'b1, 1'b0};
328: data_out = {8'd41, 8'd28, 1'b1, 1'b0};
329: data_out = {8'd50, 8'd28, 1'b1, 1'b0};
330: data_out = {8'd53, 8'd28, 1'b1, 1'b0};
331: data_out = {8'd62, 8'd28, 1'b1, 1'b0};
332: data_out = {8'd90, 8'd28, 1'b1, 1'b0};
333: data_out = {8'd95, 8'd28, 1'b1, 1'b0};
334: data_out = {8'd102, 8'd28, 1'b1, 1'b0};
335: data_out = {8'd111, 8'd28, 1'b1, 1'b0};
336: data_out = {8'd139, 8'd28, 1'b1, 1'b0};
337: data_out = {8'd148, 8'd28, 1'b1, 1'b0};
338: data_out = {8'd155, 8'd28, 1'b1, 1'b0};
339: data_out = {8'd164, 8'd28, 1'b1, 1'b0};
340: data_out = {8'd184, 8'd28, 1'b1, 1'b0};
341: data_out = {8'd193, 8'd28, 1'b1, 1'b0};
342: data_out = {8'd204, 8'd28, 1'b1, 1'b0};
343: data_out = {8'd213, 8'd28, 1'b1, 1'b0};
344: data_out = {8'd41, 8'd29, 1'b1, 1'b0};
345: data_out = {8'd50, 8'd29, 1'b1, 1'b0};
346: data_out = {8'd53, 8'd29, 1'b1, 1'b0};
347: data_out = {8'd62, 8'd29, 1'b1, 1'b0};
348: data_out = {8'd90, 8'd29, 1'b1, 1'b0};
349: data_out = {8'd95, 8'd29, 1'b1, 1'b0};
350: data_out = {8'd102, 8'd29, 1'b1, 1'b0};
351: data_out = {8'd111, 8'd29, 1'b1, 1'b0};
352: data_out = {8'd139, 8'd29, 1'b1, 1'b0};
353: data_out = {8'd148, 8'd29, 1'b1, 1'b0};
354: data_out = {8'd155, 8'd29, 1'b1, 1'b0};
355: data_out = {8'd164, 8'd29, 1'b1, 1'b0};
356: data_out = {8'd184, 8'd29, 1'b1, 1'b0};
357: data_out = {8'd193, 8'd29, 1'b1, 1'b0};
358: data_out = {8'd204, 8'd29, 1'b1, 1'b0};
359: data_out = {8'd213, 8'd29, 1'b1, 1'b0};
360: data_out = {8'd41, 8'd30, 1'b1, 1'b0};
361: data_out = {8'd50, 8'd30, 1'b1, 1'b0};
362: data_out = {8'd53, 8'd30, 1'b1, 1'b0};
363: data_out = {8'd62, 8'd30, 1'b1, 1'b0};
364: data_out = {8'd90, 8'd30, 1'b1, 1'b0};
365: data_out = {8'd95, 8'd30, 1'b1, 1'b0};
366: data_out = {8'd102, 8'd30, 1'b1, 1'b0};
367: data_out = {8'd111, 8'd30, 1'b1, 1'b0};
368: data_out = {8'd139, 8'd30, 1'b1, 1'b0};
369: data_out = {8'd148, 8'd30, 1'b1, 1'b0};
370: data_out = {8'd155, 8'd30, 1'b1, 1'b0};
371: data_out = {8'd164, 8'd30, 1'b1, 1'b0};
372: data_out = {8'd184, 8'd30, 1'b1, 1'b0};
373: data_out = {8'd193, 8'd30, 1'b1, 1'b0};
374: data_out = {8'd204, 8'd30, 1'b1, 1'b0};
375: data_out = {8'd213, 8'd30, 1'b1, 1'b0};
376: data_out = {8'd41, 8'd31, 1'b1, 1'b0};
377: data_out = {8'd50, 8'd31, 1'b1, 1'b0};
378: data_out = {8'd51, 8'd31, 1'b1, 1'b0};
379: data_out = {8'd52, 8'd31, 1'b1, 1'b0};
380: data_out = {8'd53, 8'd31, 1'b1, 1'b0};
381: data_out = {8'd62, 8'd31, 1'b1, 1'b0};
382: data_out = {8'd90, 8'd31, 1'b1, 1'b0};
383: data_out = {8'd95, 8'd31, 1'b1, 1'b0};
384: data_out = {8'd96, 8'd31, 1'b1, 1'b0};
385: data_out = {8'd97, 8'd31, 1'b1, 1'b0};
386: data_out = {8'd98, 8'd31, 1'b1, 1'b0};
387: data_out = {8'd99, 8'd31, 1'b1, 1'b0};
388: data_out = {8'd100, 8'd31, 1'b1, 1'b0};
389: data_out = {8'd101, 8'd31, 1'b1, 1'b0};
390: data_out = {8'd102, 8'd31, 1'b1, 1'b0};
391: data_out = {8'd111, 8'd31, 1'b1, 1'b0};
392: data_out = {8'd139, 8'd31, 1'b1, 1'b0};
393: data_out = {8'd148, 8'd31, 1'b1, 1'b0};
394: data_out = {8'd155, 8'd31, 1'b1, 1'b0};
395: data_out = {8'd164, 8'd31, 1'b1, 1'b0};
396: data_out = {8'd184, 8'd31, 1'b1, 1'b0};
397: data_out = {8'd193, 8'd31, 1'b1, 1'b0};
398: data_out = {8'd204, 8'd31, 1'b1, 1'b0};
399: data_out = {8'd213, 8'd31, 1'b1, 1'b0};
400: data_out = {8'd41, 8'd32, 1'b1, 1'b0};
401: data_out = {8'd62, 8'd32, 1'b1, 1'b0};
402: data_out = {8'd90, 8'd32, 1'b1, 1'b0};
403: data_out = {8'd111, 8'd32, 1'b1, 1'b0};
404: data_out = {8'd139, 8'd32, 1'b1, 1'b0};
405: data_out = {8'd148, 8'd32, 1'b1, 1'b0};
406: data_out = {8'd155, 8'd32, 1'b1, 1'b0};
407: data_out = {8'd164, 8'd32, 1'b1, 1'b0};
408: data_out = {8'd184, 8'd32, 1'b1, 1'b0};
409: data_out = {8'd193, 8'd32, 1'b1, 1'b0};
410: data_out = {8'd204, 8'd32, 1'b1, 1'b0};
411: data_out = {8'd213, 8'd32, 1'b1, 1'b0};
412: data_out = {8'd41, 8'd33, 1'b1, 1'b0};
413: data_out = {8'd62, 8'd33, 1'b1, 1'b0};
414: data_out = {8'd90, 8'd33, 1'b1, 1'b0};
415: data_out = {8'd111, 8'd33, 1'b1, 1'b0};
416: data_out = {8'd139, 8'd33, 1'b1, 1'b0};
417: data_out = {8'd148, 8'd33, 1'b1, 1'b0};
418: data_out = {8'd155, 8'd33, 1'b1, 1'b0};
419: data_out = {8'd164, 8'd33, 1'b1, 1'b0};
420: data_out = {8'd184, 8'd33, 1'b1, 1'b0};
421: data_out = {8'd193, 8'd33, 1'b1, 1'b0};
422: data_out = {8'd204, 8'd33, 1'b1, 1'b0};
423: data_out = {8'd213, 8'd33, 1'b1, 1'b0};
424: data_out = {8'd41, 8'd34, 1'b1, 1'b0};
425: data_out = {8'd62, 8'd34, 1'b1, 1'b0};
426: data_out = {8'd90, 8'd34, 1'b1, 1'b0};
427: data_out = {8'd111, 8'd34, 1'b1, 1'b0};
428: data_out = {8'd139, 8'd34, 1'b1, 1'b0};
429: data_out = {8'd148, 8'd34, 1'b1, 1'b0};
430: data_out = {8'd155, 8'd34, 1'b1, 1'b0};
431: data_out = {8'd164, 8'd34, 1'b1, 1'b0};
432: data_out = {8'd184, 8'd34, 1'b1, 1'b0};
433: data_out = {8'd193, 8'd34, 1'b1, 1'b0};
434: data_out = {8'd204, 8'd34, 1'b1, 1'b0};
435: data_out = {8'd213, 8'd34, 1'b1, 1'b0};
436: data_out = {8'd37, 8'd35, 1'b1, 1'b0};
437: data_out = {8'd38, 8'd35, 1'b1, 1'b0};
438: data_out = {8'd39, 8'd35, 1'b1, 1'b0};
439: data_out = {8'd40, 8'd35, 1'b1, 1'b0};
440: data_out = {8'd41, 8'd35, 1'b1, 1'b0};
441: data_out = {8'd46, 8'd35, 1'b1, 1'b0};
442: data_out = {8'd47, 8'd35, 1'b1, 1'b0};
443: data_out = {8'd48, 8'd35, 1'b1, 1'b0};
444: data_out = {8'd49, 8'd35, 1'b1, 1'b0};
445: data_out = {8'd50, 8'd35, 1'b1, 1'b0};
446: data_out = {8'd51, 8'd35, 1'b1, 1'b0};
447: data_out = {8'd52, 8'd35, 1'b1, 1'b0};
448: data_out = {8'd53, 8'd35, 1'b1, 1'b0};
449: data_out = {8'd62, 8'd35, 1'b1, 1'b0};
450: data_out = {8'd90, 8'd35, 1'b1, 1'b0};
451: data_out = {8'd95, 8'd35, 1'b1, 1'b0};
452: data_out = {8'd96, 8'd35, 1'b1, 1'b0};
453: data_out = {8'd97, 8'd35, 1'b1, 1'b0};
454: data_out = {8'd98, 8'd35, 1'b1, 1'b0};
455: data_out = {8'd99, 8'd35, 1'b1, 1'b0};
456: data_out = {8'd100, 8'd35, 1'b1, 1'b0};
457: data_out = {8'd101, 8'd35, 1'b1, 1'b0};
458: data_out = {8'd102, 8'd35, 1'b1, 1'b0};
459: data_out = {8'd111, 8'd35, 1'b1, 1'b0};
460: data_out = {8'd139, 8'd35, 1'b1, 1'b0};
461: data_out = {8'd148, 8'd35, 1'b1, 1'b0};
462: data_out = {8'd155, 8'd35, 1'b1, 1'b0};
463: data_out = {8'd164, 8'd35, 1'b1, 1'b0};
464: data_out = {8'd184, 8'd35, 1'b1, 1'b0};
465: data_out = {8'd193, 8'd35, 1'b1, 1'b0};
466: data_out = {8'd204, 8'd35, 1'b1, 1'b0};
467: data_out = {8'd213, 8'd35, 1'b1, 1'b0};
468: data_out = {8'd37, 8'd36, 1'b1, 1'b0};
469: data_out = {8'd46, 8'd36, 1'b1, 1'b0};
470: data_out = {8'd53, 8'd36, 1'b1, 1'b0};
471: data_out = {8'd62, 8'd36, 1'b1, 1'b0};
472: data_out = {8'd90, 8'd36, 1'b1, 1'b0};
473: data_out = {8'd95, 8'd36, 1'b1, 1'b0};
474: data_out = {8'd102, 8'd36, 1'b1, 1'b0};
475: data_out = {8'd111, 8'd36, 1'b1, 1'b0};
476: data_out = {8'd139, 8'd36, 1'b1, 1'b0};
477: data_out = {8'd148, 8'd36, 1'b1, 1'b0};
478: data_out = {8'd155, 8'd36, 1'b1, 1'b0};
479: data_out = {8'd164, 8'd36, 1'b1, 1'b0};
480: data_out = {8'd184, 8'd36, 1'b1, 1'b0};
481: data_out = {8'd193, 8'd36, 1'b1, 1'b0};
482: data_out = {8'd204, 8'd36, 1'b1, 1'b0};
483: data_out = {8'd213, 8'd36, 1'b1, 1'b0};
484: data_out = {8'd37, 8'd37, 1'b1, 1'b0};
485: data_out = {8'd46, 8'd37, 1'b1, 1'b0};
486: data_out = {8'd53, 8'd37, 1'b1, 1'b0};
487: data_out = {8'd62, 8'd37, 1'b1, 1'b0};
488: data_out = {8'd90, 8'd37, 1'b1, 1'b0};
489: data_out = {8'd95, 8'd37, 1'b1, 1'b0};
490: data_out = {8'd102, 8'd37, 1'b1, 1'b0};
491: data_out = {8'd111, 8'd37, 1'b1, 1'b0};
492: data_out = {8'd139, 8'd37, 1'b1, 1'b0};
493: data_out = {8'd148, 8'd37, 1'b1, 1'b0};
494: data_out = {8'd155, 8'd37, 1'b1, 1'b0};
495: data_out = {8'd164, 8'd37, 1'b1, 1'b0};
496: data_out = {8'd184, 8'd37, 1'b1, 1'b0};
497: data_out = {8'd193, 8'd37, 1'b1, 1'b0};
498: data_out = {8'd204, 8'd37, 1'b1, 1'b0};
499: data_out = {8'd213, 8'd37, 1'b1, 1'b0};
500: data_out = {8'd37, 8'd38, 1'b1, 1'b0};
501: data_out = {8'd46, 8'd38, 1'b1, 1'b0};
502: data_out = {8'd53, 8'd38, 1'b1, 1'b0};
503: data_out = {8'd62, 8'd38, 1'b1, 1'b0};
504: data_out = {8'd90, 8'd38, 1'b1, 1'b0};
505: data_out = {8'd95, 8'd38, 1'b1, 1'b0};
506: data_out = {8'd102, 8'd38, 1'b1, 1'b0};
507: data_out = {8'd111, 8'd38, 1'b1, 1'b0};
508: data_out = {8'd139, 8'd38, 1'b1, 1'b0};
509: data_out = {8'd148, 8'd38, 1'b1, 1'b0};
510: data_out = {8'd155, 8'd38, 1'b1, 1'b0};
511: data_out = {8'd164, 8'd38, 1'b1, 1'b0};
512: data_out = {8'd184, 8'd38, 1'b1, 1'b0};
513: data_out = {8'd193, 8'd38, 1'b1, 1'b0};
514: data_out = {8'd204, 8'd38, 1'b1, 1'b0};
515: data_out = {8'd213, 8'd38, 1'b1, 1'b0};
516: data_out = {8'd37, 8'd39, 1'b1, 1'b0};
517: data_out = {8'd46, 8'd39, 1'b1, 1'b0};
518: data_out = {8'd53, 8'd39, 1'b1, 1'b0};
519: data_out = {8'd62, 8'd39, 1'b1, 1'b0};
520: data_out = {8'd90, 8'd39, 1'b1, 1'b0};
521: data_out = {8'd91, 8'd39, 1'b1, 1'b0};
522: data_out = {8'd92, 8'd39, 1'b1, 1'b0};
523: data_out = {8'd93, 8'd39, 1'b1, 1'b0};
524: data_out = {8'd94, 8'd39, 1'b1, 1'b0};
525: data_out = {8'd95, 8'd39, 1'b1, 1'b0};
526: data_out = {8'd102, 8'd39, 1'b1, 1'b0};
527: data_out = {8'd111, 8'd39, 1'b1, 1'b0};
528: data_out = {8'd139, 8'd39, 1'b1, 1'b0};
529: data_out = {8'd148, 8'd39, 1'b1, 1'b0};
530: data_out = {8'd155, 8'd39, 1'b1, 1'b0};
531: data_out = {8'd164, 8'd39, 1'b1, 1'b0};
532: data_out = {8'd184, 8'd39, 1'b1, 1'b0};
533: data_out = {8'd193, 8'd39, 1'b1, 1'b0};
534: data_out = {8'd204, 8'd39, 1'b1, 1'b0};
535: data_out = {8'd213, 8'd39, 1'b1, 1'b0};
536: data_out = {8'd37, 8'd40, 1'b1, 1'b0};
537: data_out = {8'd46, 8'd40, 1'b1, 1'b0};
538: data_out = {8'd53, 8'd40, 1'b1, 1'b0};
539: data_out = {8'd62, 8'd40, 1'b1, 1'b0};
540: data_out = {8'd102, 8'd40, 1'b1, 1'b0};
541: data_out = {8'd111, 8'd40, 1'b1, 1'b0};
542: data_out = {8'd139, 8'd40, 1'b1, 1'b0};
543: data_out = {8'd148, 8'd40, 1'b1, 1'b0};
544: data_out = {8'd155, 8'd40, 1'b1, 1'b0};
545: data_out = {8'd164, 8'd40, 1'b1, 1'b0};
546: data_out = {8'd184, 8'd40, 1'b1, 1'b0};
547: data_out = {8'd193, 8'd40, 1'b1, 1'b0};
548: data_out = {8'd204, 8'd40, 1'b1, 1'b0};
549: data_out = {8'd213, 8'd40, 1'b1, 1'b0};
550: data_out = {8'd37, 8'd41, 1'b1, 1'b0};
551: data_out = {8'd46, 8'd41, 1'b1, 1'b0};
552: data_out = {8'd53, 8'd41, 1'b1, 1'b0};
553: data_out = {8'd62, 8'd41, 1'b1, 1'b0};
554: data_out = {8'd102, 8'd41, 1'b1, 1'b0};
555: data_out = {8'd111, 8'd41, 1'b1, 1'b0};
556: data_out = {8'd139, 8'd41, 1'b1, 1'b0};
557: data_out = {8'd148, 8'd41, 1'b1, 1'b0};
558: data_out = {8'd155, 8'd41, 1'b1, 1'b0};
559: data_out = {8'd164, 8'd41, 1'b1, 1'b0};
560: data_out = {8'd184, 8'd41, 1'b1, 1'b0};
561: data_out = {8'd193, 8'd41, 1'b1, 1'b0};
562: data_out = {8'd204, 8'd41, 1'b1, 1'b0};
563: data_out = {8'd213, 8'd41, 1'b1, 1'b0};
564: data_out = {8'd37, 8'd42, 1'b1, 1'b0};
565: data_out = {8'd46, 8'd42, 1'b1, 1'b0};
566: data_out = {8'd53, 8'd42, 1'b1, 1'b0};
567: data_out = {8'd62, 8'd42, 1'b1, 1'b0};
568: data_out = {8'd102, 8'd42, 1'b1, 1'b0};
569: data_out = {8'd111, 8'd42, 1'b1, 1'b0};
570: data_out = {8'd139, 8'd42, 1'b1, 1'b0};
571: data_out = {8'd148, 8'd42, 1'b1, 1'b0};
572: data_out = {8'd155, 8'd42, 1'b1, 1'b0};
573: data_out = {8'd164, 8'd42, 1'b1, 1'b0};
574: data_out = {8'd184, 8'd42, 1'b1, 1'b0};
575: data_out = {8'd193, 8'd42, 1'b1, 1'b0};
576: data_out = {8'd204, 8'd42, 1'b1, 1'b0};
577: data_out = {8'd213, 8'd42, 1'b1, 1'b0};
578: data_out = {8'd37, 8'd43, 1'b1, 1'b0};
579: data_out = {8'd46, 8'd43, 1'b1, 1'b0};
580: data_out = {8'd53, 8'd43, 1'b1, 1'b0};
581: data_out = {8'd62, 8'd43, 1'b1, 1'b0};
582: data_out = {8'd86, 8'd43, 1'b1, 1'b0};
583: data_out = {8'd87, 8'd43, 1'b1, 1'b0};
584: data_out = {8'd88, 8'd43, 1'b1, 1'b0};
585: data_out = {8'd89, 8'd43, 1'b1, 1'b0};
586: data_out = {8'd90, 8'd43, 1'b1, 1'b0};
587: data_out = {8'd91, 8'd43, 1'b1, 1'b0};
588: data_out = {8'd102, 8'd43, 1'b1, 1'b0};
589: data_out = {8'd111, 8'd43, 1'b1, 1'b0};
590: data_out = {8'd139, 8'd43, 1'b1, 1'b0};
591: data_out = {8'd148, 8'd43, 1'b1, 1'b0};
592: data_out = {8'd155, 8'd43, 1'b1, 1'b0};
593: data_out = {8'd164, 8'd43, 1'b1, 1'b0};
594: data_out = {8'd184, 8'd43, 1'b1, 1'b0};
595: data_out = {8'd185, 8'd43, 1'b1, 1'b0};
596: data_out = {8'd186, 8'd43, 1'b1, 1'b0};
597: data_out = {8'd187, 8'd43, 1'b1, 1'b0};
598: data_out = {8'd188, 8'd43, 1'b1, 1'b0};
599: data_out = {8'd193, 8'd43, 1'b1, 1'b0};
600: data_out = {8'd194, 8'd43, 1'b1, 1'b0};
601: data_out = {8'd195, 8'd43, 1'b1, 1'b0};
602: data_out = {8'd196, 8'd43, 1'b1, 1'b0};
603: data_out = {8'd197, 8'd43, 1'b1, 1'b0};
604: data_out = {8'd200, 8'd43, 1'b1, 1'b0};
605: data_out = {8'd201, 8'd43, 1'b1, 1'b0};
606: data_out = {8'd202, 8'd43, 1'b1, 1'b0};
607: data_out = {8'd203, 8'd43, 1'b1, 1'b0};
608: data_out = {8'd204, 8'd43, 1'b1, 1'b0};
609: data_out = {8'd209, 8'd43, 1'b1, 1'b0};
610: data_out = {8'd210, 8'd43, 1'b1, 1'b0};
611: data_out = {8'd211, 8'd43, 1'b1, 1'b0};
612: data_out = {8'd212, 8'd43, 1'b1, 1'b0};
613: data_out = {8'd213, 8'd43, 1'b1, 1'b0};
614: data_out = {8'd37, 8'd44, 1'b1, 1'b0};
615: data_out = {8'd46, 8'd44, 1'b1, 1'b0};
616: data_out = {8'd53, 8'd44, 1'b1, 1'b0};
617: data_out = {8'd62, 8'd44, 1'b1, 1'b0};
618: data_out = {8'd86, 8'd44, 1'b1, 1'b0};
619: data_out = {8'd91, 8'd44, 1'b1, 1'b0};
620: data_out = {8'd102, 8'd44, 1'b1, 1'b0};
621: data_out = {8'd111, 8'd44, 1'b1, 1'b0};
622: data_out = {8'd139, 8'd44, 1'b1, 1'b0};
623: data_out = {8'd148, 8'd44, 1'b1, 1'b0};
624: data_out = {8'd155, 8'd44, 1'b1, 1'b0};
625: data_out = {8'd164, 8'd44, 1'b1, 1'b0};
626: data_out = {8'd188, 8'd44, 1'b1, 1'b0};
627: data_out = {8'd197, 8'd44, 1'b1, 1'b0};
628: data_out = {8'd200, 8'd44, 1'b1, 1'b0};
629: data_out = {8'd209, 8'd44, 1'b1, 1'b0};
630: data_out = {8'd37, 8'd45, 1'b1, 1'b0};
631: data_out = {8'd46, 8'd45, 1'b1, 1'b0};
632: data_out = {8'd53, 8'd45, 1'b1, 1'b0};
633: data_out = {8'd62, 8'd45, 1'b1, 1'b0};
634: data_out = {8'd86, 8'd45, 1'b1, 1'b0};
635: data_out = {8'd91, 8'd45, 1'b1, 1'b0};
636: data_out = {8'd102, 8'd45, 1'b1, 1'b0};
637: data_out = {8'd111, 8'd45, 1'b1, 1'b0};
638: data_out = {8'd139, 8'd45, 1'b1, 1'b0};
639: data_out = {8'd148, 8'd45, 1'b1, 1'b0};
640: data_out = {8'd155, 8'd45, 1'b1, 1'b0};
641: data_out = {8'd164, 8'd45, 1'b1, 1'b0};
642: data_out = {8'd188, 8'd45, 1'b1, 1'b0};
643: data_out = {8'd197, 8'd45, 1'b1, 1'b0};
644: data_out = {8'd200, 8'd45, 1'b1, 1'b0};
645: data_out = {8'd209, 8'd45, 1'b1, 1'b0};
646: data_out = {8'd37, 8'd46, 1'b1, 1'b0};
647: data_out = {8'd46, 8'd46, 1'b1, 1'b0};
648: data_out = {8'd53, 8'd46, 1'b1, 1'b0};
649: data_out = {8'd62, 8'd46, 1'b1, 1'b0};
650: data_out = {8'd86, 8'd46, 1'b1, 1'b0};
651: data_out = {8'd91, 8'd46, 1'b1, 1'b0};
652: data_out = {8'd102, 8'd46, 1'b1, 1'b0};
653: data_out = {8'd111, 8'd46, 1'b1, 1'b0};
654: data_out = {8'd139, 8'd46, 1'b1, 1'b0};
655: data_out = {8'd148, 8'd46, 1'b1, 1'b0};
656: data_out = {8'd155, 8'd46, 1'b1, 1'b0};
657: data_out = {8'd164, 8'd46, 1'b1, 1'b0};
658: data_out = {8'd188, 8'd46, 1'b1, 1'b0};
659: data_out = {8'd197, 8'd46, 1'b1, 1'b0};
660: data_out = {8'd200, 8'd46, 1'b1, 1'b0};
661: data_out = {8'd209, 8'd46, 1'b1, 1'b0};
662: data_out = {8'd37, 8'd47, 1'b1, 1'b0};
663: data_out = {8'd38, 8'd47, 1'b1, 1'b0};
664: data_out = {8'd39, 8'd47, 1'b1, 1'b0};
665: data_out = {8'd40, 8'd47, 1'b1, 1'b0};
666: data_out = {8'd41, 8'd47, 1'b1, 1'b0};
667: data_out = {8'd46, 8'd47, 1'b1, 1'b0};
668: data_out = {8'd47, 8'd47, 1'b1, 1'b0};
669: data_out = {8'd48, 8'd47, 1'b1, 1'b0};
670: data_out = {8'd49, 8'd47, 1'b1, 1'b0};
671: data_out = {8'd50, 8'd47, 1'b1, 1'b0};
672: data_out = {8'd51, 8'd47, 1'b1, 1'b0};
673: data_out = {8'd52, 8'd47, 1'b1, 1'b0};
674: data_out = {8'd53, 8'd47, 1'b1, 1'b0};
675: data_out = {8'd62, 8'd47, 1'b1, 1'b0};
676: data_out = {8'd63, 8'd47, 1'b1, 1'b0};
677: data_out = {8'd64, 8'd47, 1'b1, 1'b0};
678: data_out = {8'd65, 8'd47, 1'b1, 1'b0};
679: data_out = {8'd66, 8'd47, 1'b1, 1'b0};
680: data_out = {8'd86, 8'd47, 1'b1, 1'b0};
681: data_out = {8'd91, 8'd47, 1'b1, 1'b0};
682: data_out = {8'd92, 8'd47, 1'b1, 1'b0};
683: data_out = {8'd93, 8'd47, 1'b1, 1'b0};
684: data_out = {8'd94, 8'd47, 1'b1, 1'b0};
685: data_out = {8'd95, 8'd47, 1'b1, 1'b0};
686: data_out = {8'd96, 8'd47, 1'b1, 1'b0};
687: data_out = {8'd97, 8'd47, 1'b1, 1'b0};
688: data_out = {8'd98, 8'd47, 1'b1, 1'b0};
689: data_out = {8'd99, 8'd47, 1'b1, 1'b0};
690: data_out = {8'd100, 8'd47, 1'b1, 1'b0};
691: data_out = {8'd101, 8'd47, 1'b1, 1'b0};
692: data_out = {8'd102, 8'd47, 1'b1, 1'b0};
693: data_out = {8'd111, 8'd47, 1'b1, 1'b0};
694: data_out = {8'd112, 8'd47, 1'b1, 1'b0};
695: data_out = {8'd113, 8'd47, 1'b1, 1'b0};
696: data_out = {8'd114, 8'd47, 1'b1, 1'b0};
697: data_out = {8'd115, 8'd47, 1'b1, 1'b0};
698: data_out = {8'd139, 8'd47, 1'b1, 1'b0};
699: data_out = {8'd148, 8'd47, 1'b1, 1'b0};
700: data_out = {8'd155, 8'd47, 1'b1, 1'b0};
701: data_out = {8'd164, 8'd47, 1'b1, 1'b0};
702: data_out = {8'd188, 8'd47, 1'b1, 1'b0};
703: data_out = {8'd189, 8'd47, 1'b1, 1'b0};
704: data_out = {8'd190, 8'd47, 1'b1, 1'b0};
705: data_out = {8'd191, 8'd47, 1'b1, 1'b0};
706: data_out = {8'd192, 8'd47, 1'b1, 1'b0};
707: data_out = {8'd197, 8'd47, 1'b1, 1'b0};
708: data_out = {8'd198, 8'd47, 1'b1, 1'b0};
709: data_out = {8'd199, 8'd47, 1'b1, 1'b0};
710: data_out = {8'd200, 8'd47, 1'b1, 1'b0};
711: data_out = {8'd205, 8'd47, 1'b1, 1'b0};
712: data_out = {8'd206, 8'd47, 1'b1, 1'b0};
713: data_out = {8'd207, 8'd47, 1'b1, 1'b0};
714: data_out = {8'd208, 8'd47, 1'b1, 1'b0};
715: data_out = {8'd209, 8'd47, 1'b1, 1'b0};
716: data_out = {8'd41, 8'd48, 1'b1, 1'b0};
717: data_out = {8'd66, 8'd48, 1'b1, 1'b0};
718: data_out = {8'd86, 8'd48, 1'b1, 1'b0};
719: data_out = {8'd115, 8'd48, 1'b1, 1'b0};
720: data_out = {8'd139, 8'd48, 1'b1, 1'b0};
721: data_out = {8'd148, 8'd48, 1'b1, 1'b0};
722: data_out = {8'd155, 8'd48, 1'b1, 1'b0};
723: data_out = {8'd164, 8'd48, 1'b1, 1'b0};
724: data_out = {8'd192, 8'd48, 1'b1, 1'b0};
725: data_out = {8'd205, 8'd48, 1'b1, 1'b0};
726: data_out = {8'd41, 8'd49, 1'b1, 1'b0};
727: data_out = {8'd66, 8'd49, 1'b1, 1'b0};
728: data_out = {8'd86, 8'd49, 1'b1, 1'b0};
729: data_out = {8'd115, 8'd49, 1'b1, 1'b0};
730: data_out = {8'd139, 8'd49, 1'b1, 1'b0};
731: data_out = {8'd148, 8'd49, 1'b1, 1'b0};
732: data_out = {8'd155, 8'd49, 1'b1, 1'b0};
733: data_out = {8'd164, 8'd49, 1'b1, 1'b0};
734: data_out = {8'd192, 8'd49, 1'b1, 1'b0};
735: data_out = {8'd205, 8'd49, 1'b1, 1'b0};
736: data_out = {8'd41, 8'd50, 1'b1, 1'b0};
737: data_out = {8'd66, 8'd50, 1'b1, 1'b0};
738: data_out = {8'd86, 8'd50, 1'b1, 1'b0};
739: data_out = {8'd115, 8'd50, 1'b1, 1'b0};
740: data_out = {8'd139, 8'd50, 1'b1, 1'b0};
741: data_out = {8'd148, 8'd50, 1'b1, 1'b0};
742: data_out = {8'd155, 8'd50, 1'b1, 1'b0};
743: data_out = {8'd164, 8'd50, 1'b1, 1'b0};
744: data_out = {8'd192, 8'd50, 1'b1, 1'b0};
745: data_out = {8'd205, 8'd50, 1'b1, 1'b0};
746: data_out = {8'd41, 8'd51, 1'b1, 1'b0};
747: data_out = {8'd42, 8'd51, 1'b1, 1'b0};
748: data_out = {8'd43, 8'd51, 1'b1, 1'b0};
749: data_out = {8'd44, 8'd51, 1'b1, 1'b0};
750: data_out = {8'd45, 8'd51, 1'b1, 1'b0};
751: data_out = {8'd46, 8'd51, 1'b1, 1'b0};
752: data_out = {8'd47, 8'd51, 1'b1, 1'b0};
753: data_out = {8'd48, 8'd51, 1'b1, 1'b0};
754: data_out = {8'd49, 8'd51, 1'b1, 1'b0};
755: data_out = {8'd50, 8'd51, 1'b1, 1'b0};
756: data_out = {8'd51, 8'd51, 1'b1, 1'b0};
757: data_out = {8'd52, 8'd51, 1'b1, 1'b0};
758: data_out = {8'd53, 8'd51, 1'b1, 1'b0};
759: data_out = {8'd54, 8'd51, 1'b1, 1'b0};
760: data_out = {8'd55, 8'd51, 1'b1, 1'b0};
761: data_out = {8'd56, 8'd51, 1'b1, 1'b0};
762: data_out = {8'd57, 8'd51, 1'b1, 1'b0};
763: data_out = {8'd58, 8'd51, 1'b1, 1'b0};
764: data_out = {8'd59, 8'd51, 1'b1, 1'b0};
765: data_out = {8'd60, 8'd51, 1'b1, 1'b0};
766: data_out = {8'd61, 8'd51, 1'b1, 1'b0};
767: data_out = {8'd62, 8'd51, 1'b1, 1'b0};
768: data_out = {8'd63, 8'd51, 1'b1, 1'b0};
769: data_out = {8'd64, 8'd51, 1'b1, 1'b0};
770: data_out = {8'd65, 8'd51, 1'b1, 1'b0};
771: data_out = {8'd66, 8'd51, 1'b1, 1'b0};
772: data_out = {8'd86, 8'd51, 1'b1, 1'b0};
773: data_out = {8'd87, 8'd51, 1'b1, 1'b0};
774: data_out = {8'd88, 8'd51, 1'b1, 1'b0};
775: data_out = {8'd89, 8'd51, 1'b1, 1'b0};
776: data_out = {8'd90, 8'd51, 1'b1, 1'b0};
777: data_out = {8'd91, 8'd51, 1'b1, 1'b0};
778: data_out = {8'd92, 8'd51, 1'b1, 1'b0};
779: data_out = {8'd93, 8'd51, 1'b1, 1'b0};
780: data_out = {8'd94, 8'd51, 1'b1, 1'b0};
781: data_out = {8'd95, 8'd51, 1'b1, 1'b0};
782: data_out = {8'd96, 8'd51, 1'b1, 1'b0};
783: data_out = {8'd97, 8'd51, 1'b1, 1'b0};
784: data_out = {8'd98, 8'd51, 1'b1, 1'b0};
785: data_out = {8'd99, 8'd51, 1'b1, 1'b0};
786: data_out = {8'd100, 8'd51, 1'b1, 1'b0};
787: data_out = {8'd101, 8'd51, 1'b1, 1'b0};
788: data_out = {8'd102, 8'd51, 1'b1, 1'b0};
789: data_out = {8'd103, 8'd51, 1'b1, 1'b0};
790: data_out = {8'd104, 8'd51, 1'b1, 1'b0};
791: data_out = {8'd105, 8'd51, 1'b1, 1'b0};
792: data_out = {8'd106, 8'd51, 1'b1, 1'b0};
793: data_out = {8'd107, 8'd51, 1'b1, 1'b0};
794: data_out = {8'd108, 8'd51, 1'b1, 1'b0};
795: data_out = {8'd109, 8'd51, 1'b1, 1'b0};
796: data_out = {8'd110, 8'd51, 1'b1, 1'b0};
797: data_out = {8'd111, 8'd51, 1'b1, 1'b0};
798: data_out = {8'd112, 8'd51, 1'b1, 1'b0};
799: data_out = {8'd113, 8'd51, 1'b1, 1'b0};
800: data_out = {8'd114, 8'd51, 1'b1, 1'b0};
801: data_out = {8'd115, 8'd51, 1'b1, 1'b0};
802: data_out = {8'd139, 8'd51, 1'b1, 1'b0};
803: data_out = {8'd140, 8'd51, 1'b1, 1'b0};
804: data_out = {8'd141, 8'd51, 1'b1, 1'b0};
805: data_out = {8'd142, 8'd51, 1'b1, 1'b0};
806: data_out = {8'd143, 8'd51, 1'b1, 1'b0};
807: data_out = {8'd144, 8'd51, 1'b1, 1'b0};
808: data_out = {8'd145, 8'd51, 1'b1, 1'b0};
809: data_out = {8'd146, 8'd51, 1'b1, 1'b0};
810: data_out = {8'd147, 8'd51, 1'b1, 1'b0};
811: data_out = {8'd148, 8'd51, 1'b1, 1'b0};
812: data_out = {8'd155, 8'd51, 1'b1, 1'b0};
813: data_out = {8'd156, 8'd51, 1'b1, 1'b0};
814: data_out = {8'd157, 8'd51, 1'b1, 1'b0};
815: data_out = {8'd158, 8'd51, 1'b1, 1'b0};
816: data_out = {8'd159, 8'd51, 1'b1, 1'b0};
817: data_out = {8'd160, 8'd51, 1'b1, 1'b0};
818: data_out = {8'd161, 8'd51, 1'b1, 1'b0};
819: data_out = {8'd162, 8'd51, 1'b1, 1'b0};
820: data_out = {8'd163, 8'd51, 1'b1, 1'b0};
821: data_out = {8'd164, 8'd51, 1'b1, 1'b0};
822: data_out = {8'd192, 8'd51, 1'b1, 1'b0};
823: data_out = {8'd193, 8'd51, 1'b1, 1'b0};
824: data_out = {8'd194, 8'd51, 1'b1, 1'b0};
825: data_out = {8'd195, 8'd51, 1'b1, 1'b0};
826: data_out = {8'd196, 8'd51, 1'b1, 1'b0};
827: data_out = {8'd197, 8'd51, 1'b1, 1'b0};
828: data_out = {8'd198, 8'd51, 1'b1, 1'b0};
829: data_out = {8'd199, 8'd51, 1'b1, 1'b0};
830: data_out = {8'd200, 8'd51, 1'b1, 1'b0};
831: data_out = {8'd201, 8'd51, 1'b1, 1'b0};
832: data_out = {8'd202, 8'd51, 1'b1, 1'b0};
833: data_out = {8'd203, 8'd51, 1'b1, 1'b0};
834: data_out = {8'd204, 8'd51, 1'b1, 1'b0};
835: data_out = {8'd205, 8'd51, 1'b1, 1'b0};
836: data_out = {8'd37, 8'd79, 1'b1, 1'b0};
837: data_out = {8'd38, 8'd79, 1'b1, 1'b0};
838: data_out = {8'd39, 8'd79, 1'b1, 1'b0};
839: data_out = {8'd40, 8'd79, 1'b1, 1'b0};
840: data_out = {8'd41, 8'd79, 1'b1, 1'b0};
841: data_out = {8'd42, 8'd79, 1'b1, 1'b0};
842: data_out = {8'd43, 8'd79, 1'b1, 1'b0};
843: data_out = {8'd44, 8'd79, 1'b1, 1'b0};
844: data_out = {8'd45, 8'd79, 1'b1, 1'b0};
845: data_out = {8'd46, 8'd79, 1'b1, 1'b0};
846: data_out = {8'd47, 8'd79, 1'b1, 1'b0};
847: data_out = {8'd48, 8'd79, 1'b1, 1'b0};
848: data_out = {8'd49, 8'd79, 1'b1, 1'b0};
849: data_out = {8'd50, 8'd79, 1'b1, 1'b0};
850: data_out = {8'd51, 8'd79, 1'b1, 1'b0};
851: data_out = {8'd52, 8'd79, 1'b1, 1'b0};
852: data_out = {8'd53, 8'd79, 1'b1, 1'b0};
853: data_out = {8'd54, 8'd79, 1'b1, 1'b0};
854: data_out = {8'd55, 8'd79, 1'b1, 1'b0};
855: data_out = {8'd56, 8'd79, 1'b1, 1'b0};
856: data_out = {8'd57, 8'd79, 1'b1, 1'b0};
857: data_out = {8'd58, 8'd79, 1'b1, 1'b0};
858: data_out = {8'd59, 8'd79, 1'b1, 1'b0};
859: data_out = {8'd60, 8'd79, 1'b1, 1'b0};
860: data_out = {8'd61, 8'd79, 1'b1, 1'b0};
861: data_out = {8'd62, 8'd79, 1'b1, 1'b0};
862: data_out = {8'd63, 8'd79, 1'b1, 1'b0};
863: data_out = {8'd64, 8'd79, 1'b1, 1'b0};
864: data_out = {8'd65, 8'd79, 1'b1, 1'b0};
865: data_out = {8'd66, 8'd79, 1'b1, 1'b0};
866: data_out = {8'd86, 8'd79, 1'b1, 1'b0};
867: data_out = {8'd87, 8'd79, 1'b1, 1'b0};
868: data_out = {8'd88, 8'd79, 1'b1, 1'b0};
869: data_out = {8'd89, 8'd79, 1'b1, 1'b0};
870: data_out = {8'd90, 8'd79, 1'b1, 1'b0};
871: data_out = {8'd91, 8'd79, 1'b1, 1'b0};
872: data_out = {8'd92, 8'd79, 1'b1, 1'b0};
873: data_out = {8'd93, 8'd79, 1'b1, 1'b0};
874: data_out = {8'd94, 8'd79, 1'b1, 1'b0};
875: data_out = {8'd95, 8'd79, 1'b1, 1'b0};
876: data_out = {8'd106, 8'd79, 1'b1, 1'b0};
877: data_out = {8'd107, 8'd79, 1'b1, 1'b0};
878: data_out = {8'd108, 8'd79, 1'b1, 1'b0};
879: data_out = {8'd109, 8'd79, 1'b1, 1'b0};
880: data_out = {8'd110, 8'd79, 1'b1, 1'b0};
881: data_out = {8'd111, 8'd79, 1'b1, 1'b0};
882: data_out = {8'd112, 8'd79, 1'b1, 1'b0};
883: data_out = {8'd113, 8'd79, 1'b1, 1'b0};
884: data_out = {8'd114, 8'd79, 1'b1, 1'b0};
885: data_out = {8'd115, 8'd79, 1'b1, 1'b0};
886: data_out = {8'd139, 8'd79, 1'b1, 1'b0};
887: data_out = {8'd140, 8'd79, 1'b1, 1'b0};
888: data_out = {8'd141, 8'd79, 1'b1, 1'b0};
889: data_out = {8'd142, 8'd79, 1'b1, 1'b0};
890: data_out = {8'd143, 8'd79, 1'b1, 1'b0};
891: data_out = {8'd144, 8'd79, 1'b1, 1'b0};
892: data_out = {8'd145, 8'd79, 1'b1, 1'b0};
893: data_out = {8'd146, 8'd79, 1'b1, 1'b0};
894: data_out = {8'd147, 8'd79, 1'b1, 1'b0};
895: data_out = {8'd148, 8'd79, 1'b1, 1'b0};
896: data_out = {8'd155, 8'd79, 1'b1, 1'b0};
897: data_out = {8'd156, 8'd79, 1'b1, 1'b0};
898: data_out = {8'd157, 8'd79, 1'b1, 1'b0};
899: data_out = {8'd158, 8'd79, 1'b1, 1'b0};
900: data_out = {8'd159, 8'd79, 1'b1, 1'b0};
901: data_out = {8'd160, 8'd79, 1'b1, 1'b0};
902: data_out = {8'd161, 8'd79, 1'b1, 1'b0};
903: data_out = {8'd162, 8'd79, 1'b1, 1'b0};
904: data_out = {8'd163, 8'd79, 1'b1, 1'b0};
905: data_out = {8'd164, 8'd79, 1'b1, 1'b0};
906: data_out = {8'd184, 8'd79, 1'b1, 1'b0};
907: data_out = {8'd185, 8'd79, 1'b1, 1'b0};
908: data_out = {8'd186, 8'd79, 1'b1, 1'b0};
909: data_out = {8'd187, 8'd79, 1'b1, 1'b0};
910: data_out = {8'd188, 8'd79, 1'b1, 1'b0};
911: data_out = {8'd189, 8'd79, 1'b1, 1'b0};
912: data_out = {8'd190, 8'd79, 1'b1, 1'b0};
913: data_out = {8'd191, 8'd79, 1'b1, 1'b0};
914: data_out = {8'd192, 8'd79, 1'b1, 1'b0};
915: data_out = {8'd193, 8'd79, 1'b1, 1'b0};
916: data_out = {8'd194, 8'd79, 1'b1, 1'b0};
917: data_out = {8'd195, 8'd79, 1'b1, 1'b0};
918: data_out = {8'd196, 8'd79, 1'b1, 1'b0};
919: data_out = {8'd197, 8'd79, 1'b1, 1'b0};
920: data_out = {8'd198, 8'd79, 1'b1, 1'b0};
921: data_out = {8'd199, 8'd79, 1'b1, 1'b0};
922: data_out = {8'd200, 8'd79, 1'b1, 1'b0};
923: data_out = {8'd201, 8'd79, 1'b1, 1'b0};
924: data_out = {8'd202, 8'd79, 1'b1, 1'b0};
925: data_out = {8'd203, 8'd79, 1'b1, 1'b0};
926: data_out = {8'd204, 8'd79, 1'b1, 1'b0};
927: data_out = {8'd205, 8'd79, 1'b1, 1'b0};
928: data_out = {8'd37, 8'd80, 1'b1, 1'b0};
929: data_out = {8'd66, 8'd80, 1'b1, 1'b0};
930: data_out = {8'd86, 8'd80, 1'b1, 1'b0};
931: data_out = {8'd95, 8'd80, 1'b1, 1'b0};
932: data_out = {8'd106, 8'd80, 1'b1, 1'b0};
933: data_out = {8'd115, 8'd80, 1'b1, 1'b0};
934: data_out = {8'd139, 8'd80, 1'b1, 1'b0};
935: data_out = {8'd148, 8'd80, 1'b1, 1'b0};
936: data_out = {8'd155, 8'd80, 1'b1, 1'b0};
937: data_out = {8'd164, 8'd80, 1'b1, 1'b0};
938: data_out = {8'd184, 8'd80, 1'b1, 1'b0};
939: data_out = {8'd205, 8'd80, 1'b1, 1'b0};
940: data_out = {8'd37, 8'd81, 1'b1, 1'b0};
941: data_out = {8'd66, 8'd81, 1'b1, 1'b0};
942: data_out = {8'd86, 8'd81, 1'b1, 1'b0};
943: data_out = {8'd95, 8'd81, 1'b1, 1'b0};
944: data_out = {8'd106, 8'd81, 1'b1, 1'b0};
945: data_out = {8'd115, 8'd81, 1'b1, 1'b0};
946: data_out = {8'd139, 8'd81, 1'b1, 1'b0};
947: data_out = {8'd148, 8'd81, 1'b1, 1'b0};
948: data_out = {8'd155, 8'd81, 1'b1, 1'b0};
949: data_out = {8'd164, 8'd81, 1'b1, 1'b0};
950: data_out = {8'd184, 8'd81, 1'b1, 1'b0};
951: data_out = {8'd205, 8'd81, 1'b1, 1'b0};
952: data_out = {8'd37, 8'd82, 1'b1, 1'b0};
953: data_out = {8'd66, 8'd82, 1'b1, 1'b0};
954: data_out = {8'd86, 8'd82, 1'b1, 1'b0};
955: data_out = {8'd95, 8'd82, 1'b1, 1'b0};
956: data_out = {8'd106, 8'd82, 1'b1, 1'b0};
957: data_out = {8'd115, 8'd82, 1'b1, 1'b0};
958: data_out = {8'd139, 8'd82, 1'b1, 1'b0};
959: data_out = {8'd148, 8'd82, 1'b1, 1'b0};
960: data_out = {8'd155, 8'd82, 1'b1, 1'b0};
961: data_out = {8'd164, 8'd82, 1'b1, 1'b0};
962: data_out = {8'd184, 8'd82, 1'b1, 1'b0};
963: data_out = {8'd205, 8'd82, 1'b1, 1'b0};
964: data_out = {8'd37, 8'd83, 1'b1, 1'b0};
965: data_out = {8'd42, 8'd83, 1'b1, 1'b0};
966: data_out = {8'd43, 8'd83, 1'b1, 1'b0};
967: data_out = {8'd44, 8'd83, 1'b1, 1'b0};
968: data_out = {8'd45, 8'd83, 1'b1, 1'b0};
969: data_out = {8'd46, 8'd83, 1'b1, 1'b0};
970: data_out = {8'd47, 8'd83, 1'b1, 1'b0};
971: data_out = {8'd48, 8'd83, 1'b1, 1'b0};
972: data_out = {8'd49, 8'd83, 1'b1, 1'b0};
973: data_out = {8'd50, 8'd83, 1'b1, 1'b0};
974: data_out = {8'd51, 8'd83, 1'b1, 1'b0};
975: data_out = {8'd52, 8'd83, 1'b1, 1'b0};
976: data_out = {8'd53, 8'd83, 1'b1, 1'b0};
977: data_out = {8'd62, 8'd83, 1'b1, 1'b0};
978: data_out = {8'd63, 8'd83, 1'b1, 1'b0};
979: data_out = {8'd64, 8'd83, 1'b1, 1'b0};
980: data_out = {8'd65, 8'd83, 1'b1, 1'b0};
981: data_out = {8'd66, 8'd83, 1'b1, 1'b0};
982: data_out = {8'd86, 8'd83, 1'b1, 1'b0};
983: data_out = {8'd95, 8'd83, 1'b1, 1'b0};
984: data_out = {8'd106, 8'd83, 1'b1, 1'b0};
985: data_out = {8'd115, 8'd83, 1'b1, 1'b0};
986: data_out = {8'd139, 8'd83, 1'b1, 1'b0};
987: data_out = {8'd148, 8'd83, 1'b1, 1'b0};
988: data_out = {8'd155, 8'd83, 1'b1, 1'b0};
989: data_out = {8'd164, 8'd83, 1'b1, 1'b0};
990: data_out = {8'd184, 8'd83, 1'b1, 1'b0};
991: data_out = {8'd193, 8'd83, 1'b1, 1'b0};
992: data_out = {8'd194, 8'd83, 1'b1, 1'b0};
993: data_out = {8'd195, 8'd83, 1'b1, 1'b0};
994: data_out = {8'd196, 8'd83, 1'b1, 1'b0};
995: data_out = {8'd197, 8'd83, 1'b1, 1'b0};
996: data_out = {8'd198, 8'd83, 1'b1, 1'b0};
997: data_out = {8'd199, 8'd83, 1'b1, 1'b0};
998: data_out = {8'd200, 8'd83, 1'b1, 1'b0};
999: data_out = {8'd205, 8'd83, 1'b1, 1'b0};
1000: data_out = {8'd206, 8'd83, 1'b1, 1'b0};
1001: data_out = {8'd207, 8'd83, 1'b1, 1'b0};
1002: data_out = {8'd208, 8'd83, 1'b1, 1'b0};
1003: data_out = {8'd209, 8'd83, 1'b1, 1'b0};
1004: data_out = {8'd37, 8'd84, 1'b1, 1'b0};
1005: data_out = {8'd42, 8'd84, 1'b1, 1'b0};
1006: data_out = {8'd53, 8'd84, 1'b1, 1'b0};
1007: data_out = {8'd62, 8'd84, 1'b1, 1'b0};
1008: data_out = {8'd86, 8'd84, 1'b1, 1'b0};
1009: data_out = {8'd95, 8'd84, 1'b1, 1'b0};
1010: data_out = {8'd106, 8'd84, 1'b1, 1'b0};
1011: data_out = {8'd115, 8'd84, 1'b1, 1'b0};
1012: data_out = {8'd139, 8'd84, 1'b1, 1'b0};
1013: data_out = {8'd148, 8'd84, 1'b1, 1'b0};
1014: data_out = {8'd155, 8'd84, 1'b1, 1'b0};
1015: data_out = {8'd164, 8'd84, 1'b1, 1'b0};
1016: data_out = {8'd184, 8'd84, 1'b1, 1'b0};
1017: data_out = {8'd193, 8'd84, 1'b1, 1'b0};
1018: data_out = {8'd200, 8'd84, 1'b1, 1'b0};
1019: data_out = {8'd209, 8'd84, 1'b1, 1'b0};
1020: data_out = {8'd37, 8'd85, 1'b1, 1'b0};
1021: data_out = {8'd42, 8'd85, 1'b1, 1'b0};
1022: data_out = {8'd53, 8'd85, 1'b1, 1'b0};
1023: data_out = {8'd62, 8'd85, 1'b1, 1'b0};
1024: data_out = {8'd86, 8'd85, 1'b1, 1'b0};
1025: data_out = {8'd95, 8'd85, 1'b1, 1'b0};
1026: data_out = {8'd106, 8'd85, 1'b1, 1'b0};
1027: data_out = {8'd115, 8'd85, 1'b1, 1'b0};
1028: data_out = {8'd139, 8'd85, 1'b1, 1'b0};
1029: data_out = {8'd148, 8'd85, 1'b1, 1'b0};
1030: data_out = {8'd155, 8'd85, 1'b1, 1'b0};
1031: data_out = {8'd164, 8'd85, 1'b1, 1'b0};
1032: data_out = {8'd184, 8'd85, 1'b1, 1'b0};
1033: data_out = {8'd193, 8'd85, 1'b1, 1'b0};
1034: data_out = {8'd200, 8'd85, 1'b1, 1'b0};
1035: data_out = {8'd209, 8'd85, 1'b1, 1'b0};
1036: data_out = {8'd37, 8'd86, 1'b1, 1'b0};
1037: data_out = {8'd42, 8'd86, 1'b1, 1'b0};
1038: data_out = {8'd53, 8'd86, 1'b1, 1'b0};
1039: data_out = {8'd62, 8'd86, 1'b1, 1'b0};
1040: data_out = {8'd86, 8'd86, 1'b1, 1'b0};
1041: data_out = {8'd95, 8'd86, 1'b1, 1'b0};
1042: data_out = {8'd106, 8'd86, 1'b1, 1'b0};
1043: data_out = {8'd115, 8'd86, 1'b1, 1'b0};
1044: data_out = {8'd139, 8'd86, 1'b1, 1'b0};
1045: data_out = {8'd148, 8'd86, 1'b1, 1'b0};
1046: data_out = {8'd155, 8'd86, 1'b1, 1'b0};
1047: data_out = {8'd164, 8'd86, 1'b1, 1'b0};
1048: data_out = {8'd184, 8'd86, 1'b1, 1'b0};
1049: data_out = {8'd193, 8'd86, 1'b1, 1'b0};
1050: data_out = {8'd200, 8'd86, 1'b1, 1'b0};
1051: data_out = {8'd209, 8'd86, 1'b1, 1'b0};
1052: data_out = {8'd37, 8'd87, 1'b1, 1'b0};
1053: data_out = {8'd38, 8'd87, 1'b1, 1'b0};
1054: data_out = {8'd39, 8'd87, 1'b1, 1'b0};
1055: data_out = {8'd40, 8'd87, 1'b1, 1'b0};
1056: data_out = {8'd41, 8'd87, 1'b1, 1'b0};
1057: data_out = {8'd42, 8'd87, 1'b1, 1'b0};
1058: data_out = {8'd53, 8'd87, 1'b1, 1'b0};
1059: data_out = {8'd62, 8'd87, 1'b1, 1'b0};
1060: data_out = {8'd86, 8'd87, 1'b1, 1'b0};
1061: data_out = {8'd95, 8'd87, 1'b1, 1'b0};
1062: data_out = {8'd106, 8'd87, 1'b1, 1'b0};
1063: data_out = {8'd115, 8'd87, 1'b1, 1'b0};
1064: data_out = {8'd139, 8'd87, 1'b1, 1'b0};
1065: data_out = {8'd148, 8'd87, 1'b1, 1'b0};
1066: data_out = {8'd155, 8'd87, 1'b1, 1'b0};
1067: data_out = {8'd164, 8'd87, 1'b1, 1'b0};
1068: data_out = {8'd184, 8'd87, 1'b1, 1'b0};
1069: data_out = {8'd193, 8'd87, 1'b1, 1'b0};
1070: data_out = {8'd200, 8'd87, 1'b1, 1'b0};
1071: data_out = {8'd201, 8'd87, 1'b1, 1'b0};
1072: data_out = {8'd202, 8'd87, 1'b1, 1'b0};
1073: data_out = {8'd203, 8'd87, 1'b1, 1'b0};
1074: data_out = {8'd204, 8'd87, 1'b1, 1'b0};
1075: data_out = {8'd209, 8'd87, 1'b1, 1'b0};
1076: data_out = {8'd210, 8'd87, 1'b1, 1'b0};
1077: data_out = {8'd211, 8'd87, 1'b1, 1'b0};
1078: data_out = {8'd212, 8'd87, 1'b1, 1'b0};
1079: data_out = {8'd213, 8'd87, 1'b1, 1'b0};
1080: data_out = {8'd53, 8'd88, 1'b1, 1'b0};
1081: data_out = {8'd62, 8'd88, 1'b1, 1'b0};
1082: data_out = {8'd86, 8'd88, 1'b1, 1'b0};
1083: data_out = {8'd95, 8'd88, 1'b1, 1'b0};
1084: data_out = {8'd106, 8'd88, 1'b1, 1'b0};
1085: data_out = {8'd115, 8'd88, 1'b1, 1'b0};
1086: data_out = {8'd139, 8'd88, 1'b1, 1'b0};
1087: data_out = {8'd148, 8'd88, 1'b1, 1'b0};
1088: data_out = {8'd155, 8'd88, 1'b1, 1'b0};
1089: data_out = {8'd164, 8'd88, 1'b1, 1'b0};
1090: data_out = {8'd184, 8'd88, 1'b1, 1'b0};
1091: data_out = {8'd193, 8'd88, 1'b1, 1'b0};
1092: data_out = {8'd204, 8'd88, 1'b1, 1'b0};
1093: data_out = {8'd213, 8'd88, 1'b1, 1'b0};
1094: data_out = {8'd53, 8'd89, 1'b1, 1'b0};
1095: data_out = {8'd62, 8'd89, 1'b1, 1'b0};
1096: data_out = {8'd86, 8'd89, 1'b1, 1'b0};
1097: data_out = {8'd95, 8'd89, 1'b1, 1'b0};
1098: data_out = {8'd106, 8'd89, 1'b1, 1'b0};
1099: data_out = {8'd115, 8'd89, 1'b1, 1'b0};
1100: data_out = {8'd139, 8'd89, 1'b1, 1'b0};
1101: data_out = {8'd148, 8'd89, 1'b1, 1'b0};
1102: data_out = {8'd155, 8'd89, 1'b1, 1'b0};
1103: data_out = {8'd164, 8'd89, 1'b1, 1'b0};
1104: data_out = {8'd184, 8'd89, 1'b1, 1'b0};
1105: data_out = {8'd193, 8'd89, 1'b1, 1'b0};
1106: data_out = {8'd204, 8'd89, 1'b1, 1'b0};
1107: data_out = {8'd213, 8'd89, 1'b1, 1'b0};
1108: data_out = {8'd53, 8'd90, 1'b1, 1'b0};
1109: data_out = {8'd62, 8'd90, 1'b1, 1'b0};
1110: data_out = {8'd86, 8'd90, 1'b1, 1'b0};
1111: data_out = {8'd95, 8'd90, 1'b1, 1'b0};
1112: data_out = {8'd106, 8'd90, 1'b1, 1'b0};
1113: data_out = {8'd115, 8'd90, 1'b1, 1'b0};
1114: data_out = {8'd139, 8'd90, 1'b1, 1'b0};
1115: data_out = {8'd148, 8'd90, 1'b1, 1'b0};
1116: data_out = {8'd155, 8'd90, 1'b1, 1'b0};
1117: data_out = {8'd164, 8'd90, 1'b1, 1'b0};
1118: data_out = {8'd184, 8'd90, 1'b1, 1'b0};
1119: data_out = {8'd193, 8'd90, 1'b1, 1'b0};
1120: data_out = {8'd204, 8'd90, 1'b1, 1'b0};
1121: data_out = {8'd213, 8'd90, 1'b1, 1'b0};
1122: data_out = {8'd41, 8'd91, 1'b1, 1'b0};
1123: data_out = {8'd42, 8'd91, 1'b1, 1'b0};
1124: data_out = {8'd43, 8'd91, 1'b1, 1'b0};
1125: data_out = {8'd44, 8'd91, 1'b1, 1'b0};
1126: data_out = {8'd45, 8'd91, 1'b1, 1'b0};
1127: data_out = {8'd46, 8'd91, 1'b1, 1'b0};
1128: data_out = {8'd53, 8'd91, 1'b1, 1'b0};
1129: data_out = {8'd62, 8'd91, 1'b1, 1'b0};
1130: data_out = {8'd86, 8'd91, 1'b1, 1'b0};
1131: data_out = {8'd95, 8'd91, 1'b1, 1'b0};
1132: data_out = {8'd106, 8'd91, 1'b1, 1'b0};
1133: data_out = {8'd115, 8'd91, 1'b1, 1'b0};
1134: data_out = {8'd139, 8'd91, 1'b1, 1'b0};
1135: data_out = {8'd148, 8'd91, 1'b1, 1'b0};
1136: data_out = {8'd149, 8'd91, 1'b1, 1'b0};
1137: data_out = {8'd150, 8'd91, 1'b1, 1'b0};
1138: data_out = {8'd151, 8'd91, 1'b1, 1'b0};
1139: data_out = {8'd152, 8'd91, 1'b1, 1'b0};
1140: data_out = {8'd153, 8'd91, 1'b1, 1'b0};
1141: data_out = {8'd154, 8'd91, 1'b1, 1'b0};
1142: data_out = {8'd155, 8'd91, 1'b1, 1'b0};
1143: data_out = {8'd164, 8'd91, 1'b1, 1'b0};
1144: data_out = {8'd184, 8'd91, 1'b1, 1'b0};
1145: data_out = {8'd193, 8'd91, 1'b1, 1'b0};
1146: data_out = {8'd194, 8'd91, 1'b1, 1'b0};
1147: data_out = {8'd195, 8'd91, 1'b1, 1'b0};
1148: data_out = {8'd196, 8'd91, 1'b1, 1'b0};
1149: data_out = {8'd197, 8'd91, 1'b1, 1'b0};
1150: data_out = {8'd204, 8'd91, 1'b1, 1'b0};
1151: data_out = {8'd213, 8'd91, 1'b1, 1'b0};
1152: data_out = {8'd41, 8'd92, 1'b1, 1'b0};
1153: data_out = {8'd46, 8'd92, 1'b1, 1'b0};
1154: data_out = {8'd53, 8'd92, 1'b1, 1'b0};
1155: data_out = {8'd62, 8'd92, 1'b1, 1'b0};
1156: data_out = {8'd86, 8'd92, 1'b1, 1'b0};
1157: data_out = {8'd95, 8'd92, 1'b1, 1'b0};
1158: data_out = {8'd106, 8'd92, 1'b1, 1'b0};
1159: data_out = {8'd115, 8'd92, 1'b1, 1'b0};
1160: data_out = {8'd139, 8'd92, 1'b1, 1'b0};
1161: data_out = {8'd164, 8'd92, 1'b1, 1'b0};
1162: data_out = {8'd184, 8'd92, 1'b1, 1'b0};
1163: data_out = {8'd197, 8'd92, 1'b1, 1'b0};
1164: data_out = {8'd204, 8'd92, 1'b1, 1'b0};
1165: data_out = {8'd213, 8'd92, 1'b1, 1'b0};
1166: data_out = {8'd41, 8'd93, 1'b1, 1'b0};
1167: data_out = {8'd46, 8'd93, 1'b1, 1'b0};
1168: data_out = {8'd53, 8'd93, 1'b1, 1'b0};
1169: data_out = {8'd62, 8'd93, 1'b1, 1'b0};
1170: data_out = {8'd86, 8'd93, 1'b1, 1'b0};
1171: data_out = {8'd95, 8'd93, 1'b1, 1'b0};
1172: data_out = {8'd106, 8'd93, 1'b1, 1'b0};
1173: data_out = {8'd115, 8'd93, 1'b1, 1'b0};
1174: data_out = {8'd139, 8'd93, 1'b1, 1'b0};
1175: data_out = {8'd164, 8'd93, 1'b1, 1'b0};
1176: data_out = {8'd184, 8'd93, 1'b1, 1'b0};
1177: data_out = {8'd197, 8'd93, 1'b1, 1'b0};
1178: data_out = {8'd204, 8'd93, 1'b1, 1'b0};
1179: data_out = {8'd213, 8'd93, 1'b1, 1'b0};
1180: data_out = {8'd41, 8'd94, 1'b1, 1'b0};
1181: data_out = {8'd46, 8'd94, 1'b1, 1'b0};
1182: data_out = {8'd53, 8'd94, 1'b1, 1'b0};
1183: data_out = {8'd62, 8'd94, 1'b1, 1'b0};
1184: data_out = {8'd86, 8'd94, 1'b1, 1'b0};
1185: data_out = {8'd95, 8'd94, 1'b1, 1'b0};
1186: data_out = {8'd106, 8'd94, 1'b1, 1'b0};
1187: data_out = {8'd115, 8'd94, 1'b1, 1'b0};
1188: data_out = {8'd139, 8'd94, 1'b1, 1'b0};
1189: data_out = {8'd164, 8'd94, 1'b1, 1'b0};
1190: data_out = {8'd184, 8'd94, 1'b1, 1'b0};
1191: data_out = {8'd197, 8'd94, 1'b1, 1'b0};
1192: data_out = {8'd204, 8'd94, 1'b1, 1'b0};
1193: data_out = {8'd213, 8'd94, 1'b1, 1'b0};
1194: data_out = {8'd41, 8'd95, 1'b1, 1'b0};
1195: data_out = {8'd46, 8'd95, 1'b1, 1'b0};
1196: data_out = {8'd47, 8'd95, 1'b1, 1'b0};
1197: data_out = {8'd48, 8'd95, 1'b1, 1'b0};
1198: data_out = {8'd49, 8'd95, 1'b1, 1'b0};
1199: data_out = {8'd50, 8'd95, 1'b1, 1'b0};
1200: data_out = {8'd51, 8'd95, 1'b1, 1'b0};
1201: data_out = {8'd52, 8'd95, 1'b1, 1'b0};
1202: data_out = {8'd53, 8'd95, 1'b1, 1'b0};
1203: data_out = {8'd62, 8'd95, 1'b1, 1'b0};
1204: data_out = {8'd86, 8'd95, 1'b1, 1'b0};
1205: data_out = {8'd95, 8'd95, 1'b1, 1'b0};
1206: data_out = {8'd98, 8'd95, 1'b1, 1'b0};
1207: data_out = {8'd99, 8'd95, 1'b1, 1'b0};
1208: data_out = {8'd100, 8'd95, 1'b1, 1'b0};
1209: data_out = {8'd101, 8'd95, 1'b1, 1'b0};
1210: data_out = {8'd102, 8'd95, 1'b1, 1'b0};
1211: data_out = {8'd103, 8'd95, 1'b1, 1'b0};
1212: data_out = {8'd106, 8'd95, 1'b1, 1'b0};
1213: data_out = {8'd115, 8'd95, 1'b1, 1'b0};
1214: data_out = {8'd139, 8'd95, 1'b1, 1'b0};
1215: data_out = {8'd148, 8'd95, 1'b1, 1'b0};
1216: data_out = {8'd149, 8'd95, 1'b1, 1'b0};
1217: data_out = {8'd150, 8'd95, 1'b1, 1'b0};
1218: data_out = {8'd151, 8'd95, 1'b1, 1'b0};
1219: data_out = {8'd152, 8'd95, 1'b1, 1'b0};
1220: data_out = {8'd153, 8'd95, 1'b1, 1'b0};
1221: data_out = {8'd154, 8'd95, 1'b1, 1'b0};
1222: data_out = {8'd155, 8'd95, 1'b1, 1'b0};
1223: data_out = {8'd164, 8'd95, 1'b1, 1'b0};
1224: data_out = {8'd184, 8'd95, 1'b1, 1'b0};
1225: data_out = {8'd185, 8'd95, 1'b1, 1'b0};
1226: data_out = {8'd186, 8'd95, 1'b1, 1'b0};
1227: data_out = {8'd187, 8'd95, 1'b1, 1'b0};
1228: data_out = {8'd188, 8'd95, 1'b1, 1'b0};
1229: data_out = {8'd189, 8'd95, 1'b1, 1'b0};
1230: data_out = {8'd190, 8'd95, 1'b1, 1'b0};
1231: data_out = {8'd191, 8'd95, 1'b1, 1'b0};
1232: data_out = {8'd192, 8'd95, 1'b1, 1'b0};
1233: data_out = {8'd193, 8'd95, 1'b1, 1'b0};
1234: data_out = {8'd194, 8'd95, 1'b1, 1'b0};
1235: data_out = {8'd195, 8'd95, 1'b1, 1'b0};
1236: data_out = {8'd196, 8'd95, 1'b1, 1'b0};
1237: data_out = {8'd197, 8'd95, 1'b1, 1'b0};
1238: data_out = {8'd204, 8'd95, 1'b1, 1'b0};
1239: data_out = {8'd213, 8'd95, 1'b1, 1'b0};
1240: data_out = {8'd41, 8'd96, 1'b1, 1'b0};
1241: data_out = {8'd62, 8'd96, 1'b1, 1'b0};
1242: data_out = {8'd86, 8'd96, 1'b1, 1'b0};
1243: data_out = {8'd95, 8'd96, 1'b1, 1'b0};
1244: data_out = {8'd98, 8'd96, 1'b1, 1'b0};
1245: data_out = {8'd103, 8'd96, 1'b1, 1'b0};
1246: data_out = {8'd106, 8'd96, 1'b1, 1'b0};
1247: data_out = {8'd115, 8'd96, 1'b1, 1'b0};
1248: data_out = {8'd139, 8'd96, 1'b1, 1'b0};
1249: data_out = {8'd148, 8'd96, 1'b1, 1'b0};
1250: data_out = {8'd155, 8'd96, 1'b1, 1'b0};
1251: data_out = {8'd164, 8'd96, 1'b1, 1'b0};
1252: data_out = {8'd204, 8'd96, 1'b1, 1'b0};
1253: data_out = {8'd213, 8'd96, 1'b1, 1'b0};
1254: data_out = {8'd41, 8'd97, 1'b1, 1'b0};
1255: data_out = {8'd62, 8'd97, 1'b1, 1'b0};
1256: data_out = {8'd86, 8'd97, 1'b1, 1'b0};
1257: data_out = {8'd95, 8'd97, 1'b1, 1'b0};
1258: data_out = {8'd98, 8'd97, 1'b1, 1'b0};
1259: data_out = {8'd103, 8'd97, 1'b1, 1'b0};
1260: data_out = {8'd106, 8'd97, 1'b1, 1'b0};
1261: data_out = {8'd115, 8'd97, 1'b1, 1'b0};
1262: data_out = {8'd139, 8'd97, 1'b1, 1'b0};
1263: data_out = {8'd148, 8'd97, 1'b1, 1'b0};
1264: data_out = {8'd155, 8'd97, 1'b1, 1'b0};
1265: data_out = {8'd164, 8'd97, 1'b1, 1'b0};
1266: data_out = {8'd204, 8'd97, 1'b1, 1'b0};
1267: data_out = {8'd213, 8'd97, 1'b1, 1'b0};
1268: data_out = {8'd41, 8'd98, 1'b1, 1'b0};
1269: data_out = {8'd62, 8'd98, 1'b1, 1'b0};
1270: data_out = {8'd86, 8'd98, 1'b1, 1'b0};
1271: data_out = {8'd95, 8'd98, 1'b1, 1'b0};
1272: data_out = {8'd98, 8'd98, 1'b1, 1'b0};
1273: data_out = {8'd103, 8'd98, 1'b1, 1'b0};
1274: data_out = {8'd106, 8'd98, 1'b1, 1'b0};
1275: data_out = {8'd115, 8'd98, 1'b1, 1'b0};
1276: data_out = {8'd139, 8'd98, 1'b1, 1'b0};
1277: data_out = {8'd148, 8'd98, 1'b1, 1'b0};
1278: data_out = {8'd155, 8'd98, 1'b1, 1'b0};
1279: data_out = {8'd164, 8'd98, 1'b1, 1'b0};
1280: data_out = {8'd204, 8'd98, 1'b1, 1'b0};
1281: data_out = {8'd213, 8'd98, 1'b1, 1'b0};
1282: data_out = {8'd41, 8'd99, 1'b1, 1'b0};
1283: data_out = {8'd46, 8'd99, 1'b1, 1'b0};
1284: data_out = {8'd47, 8'd99, 1'b1, 1'b0};
1285: data_out = {8'd48, 8'd99, 1'b1, 1'b0};
1286: data_out = {8'd49, 8'd99, 1'b1, 1'b0};
1287: data_out = {8'd50, 8'd99, 1'b1, 1'b0};
1288: data_out = {8'd51, 8'd99, 1'b1, 1'b0};
1289: data_out = {8'd52, 8'd99, 1'b1, 1'b0};
1290: data_out = {8'd53, 8'd99, 1'b1, 1'b0};
1291: data_out = {8'd62, 8'd99, 1'b1, 1'b0};
1292: data_out = {8'd86, 8'd99, 1'b1, 1'b0};
1293: data_out = {8'd95, 8'd99, 1'b1, 1'b0};
1294: data_out = {8'd96, 8'd99, 1'b1, 1'b0};
1295: data_out = {8'd97, 8'd99, 1'b1, 1'b0};
1296: data_out = {8'd98, 8'd99, 1'b1, 1'b0};
1297: data_out = {8'd103, 8'd99, 1'b1, 1'b0};
1298: data_out = {8'd104, 8'd99, 1'b1, 1'b0};
1299: data_out = {8'd105, 8'd99, 1'b1, 1'b0};
1300: data_out = {8'd106, 8'd99, 1'b1, 1'b0};
1301: data_out = {8'd115, 8'd99, 1'b1, 1'b0};
1302: data_out = {8'd139, 8'd99, 1'b1, 1'b0};
1303: data_out = {8'd148, 8'd99, 1'b1, 1'b0};
1304: data_out = {8'd155, 8'd99, 1'b1, 1'b0};
1305: data_out = {8'd164, 8'd99, 1'b1, 1'b0};
1306: data_out = {8'd204, 8'd99, 1'b1, 1'b0};
1307: data_out = {8'd213, 8'd99, 1'b1, 1'b0};
1308: data_out = {8'd41, 8'd100, 1'b1, 1'b0};
1309: data_out = {8'd46, 8'd100, 1'b1, 1'b0};
1310: data_out = {8'd53, 8'd100, 1'b1, 1'b0};
1311: data_out = {8'd62, 8'd100, 1'b1, 1'b0};
1312: data_out = {8'd86, 8'd100, 1'b1, 1'b0};
1313: data_out = {8'd115, 8'd100, 1'b1, 1'b0};
1314: data_out = {8'd139, 8'd100, 1'b1, 1'b0};
1315: data_out = {8'd148, 8'd100, 1'b1, 1'b0};
1316: data_out = {8'd155, 8'd100, 1'b1, 1'b0};
1317: data_out = {8'd164, 8'd100, 1'b1, 1'b0};
1318: data_out = {8'd204, 8'd100, 1'b1, 1'b0};
1319: data_out = {8'd213, 8'd100, 1'b1, 1'b0};
1320: data_out = {8'd41, 8'd101, 1'b1, 1'b0};
1321: data_out = {8'd46, 8'd101, 1'b1, 1'b0};
1322: data_out = {8'd53, 8'd101, 1'b1, 1'b0};
1323: data_out = {8'd62, 8'd101, 1'b1, 1'b0};
1324: data_out = {8'd86, 8'd101, 1'b1, 1'b0};
1325: data_out = {8'd115, 8'd101, 1'b1, 1'b0};
1326: data_out = {8'd139, 8'd101, 1'b1, 1'b0};
1327: data_out = {8'd148, 8'd101, 1'b1, 1'b0};
1328: data_out = {8'd155, 8'd101, 1'b1, 1'b0};
1329: data_out = {8'd164, 8'd101, 1'b1, 1'b0};
1330: data_out = {8'd204, 8'd101, 1'b1, 1'b0};
1331: data_out = {8'd213, 8'd101, 1'b1, 1'b0};
1332: data_out = {8'd41, 8'd102, 1'b1, 1'b0};
1333: data_out = {8'd46, 8'd102, 1'b1, 1'b0};
1334: data_out = {8'd53, 8'd102, 1'b1, 1'b0};
1335: data_out = {8'd62, 8'd102, 1'b1, 1'b0};
1336: data_out = {8'd86, 8'd102, 1'b1, 1'b0};
1337: data_out = {8'd115, 8'd102, 1'b1, 1'b0};
1338: data_out = {8'd139, 8'd102, 1'b1, 1'b0};
1339: data_out = {8'd148, 8'd102, 1'b1, 1'b0};
1340: data_out = {8'd155, 8'd102, 1'b1, 1'b0};
1341: data_out = {8'd164, 8'd102, 1'b1, 1'b0};
1342: data_out = {8'd204, 8'd102, 1'b1, 1'b0};
1343: data_out = {8'd213, 8'd102, 1'b1, 1'b0};
1344: data_out = {8'd41, 8'd103, 1'b1, 1'b0};
1345: data_out = {8'd42, 8'd103, 1'b1, 1'b0};
1346: data_out = {8'd43, 8'd103, 1'b1, 1'b0};
1347: data_out = {8'd44, 8'd103, 1'b1, 1'b0};
1348: data_out = {8'd45, 8'd103, 1'b1, 1'b0};
1349: data_out = {8'd46, 8'd103, 1'b1, 1'b0};
1350: data_out = {8'd53, 8'd103, 1'b1, 1'b0};
1351: data_out = {8'd62, 8'd103, 1'b1, 1'b0};
1352: data_out = {8'd86, 8'd103, 1'b1, 1'b0};
1353: data_out = {8'd115, 8'd103, 1'b1, 1'b0};
1354: data_out = {8'd139, 8'd103, 1'b1, 1'b0};
1355: data_out = {8'd148, 8'd103, 1'b1, 1'b0};
1356: data_out = {8'd155, 8'd103, 1'b1, 1'b0};
1357: data_out = {8'd164, 8'd103, 1'b1, 1'b0};
1358: data_out = {8'd184, 8'd103, 1'b1, 1'b0};
1359: data_out = {8'd185, 8'd103, 1'b1, 1'b0};
1360: data_out = {8'd186, 8'd103, 1'b1, 1'b0};
1361: data_out = {8'd187, 8'd103, 1'b1, 1'b0};
1362: data_out = {8'd188, 8'd103, 1'b1, 1'b0};
1363: data_out = {8'd189, 8'd103, 1'b1, 1'b0};
1364: data_out = {8'd190, 8'd103, 1'b1, 1'b0};
1365: data_out = {8'd191, 8'd103, 1'b1, 1'b0};
1366: data_out = {8'd192, 8'd103, 1'b1, 1'b0};
1367: data_out = {8'd193, 8'd103, 1'b1, 1'b0};
1368: data_out = {8'd204, 8'd103, 1'b1, 1'b0};
1369: data_out = {8'd213, 8'd103, 1'b1, 1'b0};
1370: data_out = {8'd53, 8'd104, 1'b1, 1'b0};
1371: data_out = {8'd62, 8'd104, 1'b1, 1'b0};
1372: data_out = {8'd86, 8'd104, 1'b1, 1'b0};
1373: data_out = {8'd115, 8'd104, 1'b1, 1'b0};
1374: data_out = {8'd139, 8'd104, 1'b1, 1'b0};
1375: data_out = {8'd148, 8'd104, 1'b1, 1'b0};
1376: data_out = {8'd155, 8'd104, 1'b1, 1'b0};
1377: data_out = {8'd164, 8'd104, 1'b1, 1'b0};
1378: data_out = {8'd184, 8'd104, 1'b1, 1'b0};
1379: data_out = {8'd193, 8'd104, 1'b1, 1'b0};
1380: data_out = {8'd204, 8'd104, 1'b1, 1'b0};
1381: data_out = {8'd213, 8'd104, 1'b1, 1'b0};
1382: data_out = {8'd53, 8'd105, 1'b1, 1'b0};
1383: data_out = {8'd62, 8'd105, 1'b1, 1'b0};
1384: data_out = {8'd86, 8'd105, 1'b1, 1'b0};
1385: data_out = {8'd115, 8'd105, 1'b1, 1'b0};
1386: data_out = {8'd139, 8'd105, 1'b1, 1'b0};
1387: data_out = {8'd148, 8'd105, 1'b1, 1'b0};
1388: data_out = {8'd155, 8'd105, 1'b1, 1'b0};
1389: data_out = {8'd164, 8'd105, 1'b1, 1'b0};
1390: data_out = {8'd184, 8'd105, 1'b1, 1'b0};
1391: data_out = {8'd193, 8'd105, 1'b1, 1'b0};
1392: data_out = {8'd204, 8'd105, 1'b1, 1'b0};
1393: data_out = {8'd213, 8'd105, 1'b1, 1'b0};
1394: data_out = {8'd53, 8'd106, 1'b1, 1'b0};
1395: data_out = {8'd62, 8'd106, 1'b1, 1'b0};
1396: data_out = {8'd86, 8'd106, 1'b1, 1'b0};
1397: data_out = {8'd115, 8'd106, 1'b1, 1'b0};
1398: data_out = {8'd139, 8'd106, 1'b1, 1'b0};
1399: data_out = {8'd148, 8'd106, 1'b1, 1'b0};
1400: data_out = {8'd155, 8'd106, 1'b1, 1'b0};
1401: data_out = {8'd164, 8'd106, 1'b1, 1'b0};
1402: data_out = {8'd184, 8'd106, 1'b1, 1'b0};
1403: data_out = {8'd193, 8'd106, 1'b1, 1'b0};
1404: data_out = {8'd204, 8'd106, 1'b1, 1'b0};
1405: data_out = {8'd213, 8'd106, 1'b1, 1'b0};
1406: data_out = {8'd37, 8'd107, 1'b1, 1'b0};
1407: data_out = {8'd38, 8'd107, 1'b1, 1'b0};
1408: data_out = {8'd39, 8'd107, 1'b1, 1'b0};
1409: data_out = {8'd40, 8'd107, 1'b1, 1'b0};
1410: data_out = {8'd41, 8'd107, 1'b1, 1'b0};
1411: data_out = {8'd42, 8'd107, 1'b1, 1'b0};
1412: data_out = {8'd53, 8'd107, 1'b1, 1'b0};
1413: data_out = {8'd62, 8'd107, 1'b1, 1'b0};
1414: data_out = {8'd86, 8'd107, 1'b1, 1'b0};
1415: data_out = {8'd99, 8'd107, 1'b1, 1'b0};
1416: data_out = {8'd100, 8'd107, 1'b1, 1'b0};
1417: data_out = {8'd101, 8'd107, 1'b1, 1'b0};
1418: data_out = {8'd102, 8'd107, 1'b1, 1'b0};
1419: data_out = {8'd115, 8'd107, 1'b1, 1'b0};
1420: data_out = {8'd139, 8'd107, 1'b1, 1'b0};
1421: data_out = {8'd140, 8'd107, 1'b1, 1'b0};
1422: data_out = {8'd141, 8'd107, 1'b1, 1'b0};
1423: data_out = {8'd142, 8'd107, 1'b1, 1'b0};
1424: data_out = {8'd143, 8'd107, 1'b1, 1'b0};
1425: data_out = {8'd148, 8'd107, 1'b1, 1'b0};
1426: data_out = {8'd149, 8'd107, 1'b1, 1'b0};
1427: data_out = {8'd150, 8'd107, 1'b1, 1'b0};
1428: data_out = {8'd151, 8'd107, 1'b1, 1'b0};
1429: data_out = {8'd152, 8'd107, 1'b1, 1'b0};
1430: data_out = {8'd153, 8'd107, 1'b1, 1'b0};
1431: data_out = {8'd154, 8'd107, 1'b1, 1'b0};
1432: data_out = {8'd155, 8'd107, 1'b1, 1'b0};
1433: data_out = {8'd160, 8'd107, 1'b1, 1'b0};
1434: data_out = {8'd161, 8'd107, 1'b1, 1'b0};
1435: data_out = {8'd162, 8'd107, 1'b1, 1'b0};
1436: data_out = {8'd163, 8'd107, 1'b1, 1'b0};
1437: data_out = {8'd164, 8'd107, 1'b1, 1'b0};
1438: data_out = {8'd184, 8'd107, 1'b1, 1'b0};
1439: data_out = {8'd193, 8'd107, 1'b1, 1'b0};
1440: data_out = {8'd200, 8'd107, 1'b1, 1'b0};
1441: data_out = {8'd201, 8'd107, 1'b1, 1'b0};
1442: data_out = {8'd202, 8'd107, 1'b1, 1'b0};
1443: data_out = {8'd203, 8'd107, 1'b1, 1'b0};
1444: data_out = {8'd204, 8'd107, 1'b1, 1'b0};
1445: data_out = {8'd209, 8'd107, 1'b1, 1'b0};
1446: data_out = {8'd210, 8'd107, 1'b1, 1'b0};
1447: data_out = {8'd211, 8'd107, 1'b1, 1'b0};
1448: data_out = {8'd212, 8'd107, 1'b1, 1'b0};
1449: data_out = {8'd213, 8'd107, 1'b1, 1'b0};
1450: data_out = {8'd37, 8'd108, 1'b1, 1'b0};
1451: data_out = {8'd42, 8'd108, 1'b1, 1'b0};
1452: data_out = {8'd53, 8'd108, 1'b1, 1'b0};
1453: data_out = {8'd62, 8'd108, 1'b1, 1'b0};
1454: data_out = {8'd86, 8'd108, 1'b1, 1'b0};
1455: data_out = {8'd99, 8'd108, 1'b1, 1'b0};
1456: data_out = {8'd102, 8'd108, 1'b1, 1'b0};
1457: data_out = {8'd115, 8'd108, 1'b1, 1'b0};
1458: data_out = {8'd143, 8'd108, 1'b1, 1'b0};
1459: data_out = {8'd160, 8'd108, 1'b1, 1'b0};
1460: data_out = {8'd184, 8'd108, 1'b1, 1'b0};
1461: data_out = {8'd193, 8'd108, 1'b1, 1'b0};
1462: data_out = {8'd200, 8'd108, 1'b1, 1'b0};
1463: data_out = {8'd209, 8'd108, 1'b1, 1'b0};
1464: data_out = {8'd37, 8'd109, 1'b1, 1'b0};
1465: data_out = {8'd42, 8'd109, 1'b1, 1'b0};
1466: data_out = {8'd53, 8'd109, 1'b1, 1'b0};
1467: data_out = {8'd62, 8'd109, 1'b1, 1'b0};
1468: data_out = {8'd86, 8'd109, 1'b1, 1'b0};
1469: data_out = {8'd99, 8'd109, 1'b1, 1'b0};
1470: data_out = {8'd102, 8'd109, 1'b1, 1'b0};
1471: data_out = {8'd115, 8'd109, 1'b1, 1'b0};
1472: data_out = {8'd143, 8'd109, 1'b1, 1'b0};
1473: data_out = {8'd160, 8'd109, 1'b1, 1'b0};
1474: data_out = {8'd184, 8'd109, 1'b1, 1'b0};
1475: data_out = {8'd193, 8'd109, 1'b1, 1'b0};
1476: data_out = {8'd200, 8'd109, 1'b1, 1'b0};
1477: data_out = {8'd209, 8'd109, 1'b1, 1'b0};
1478: data_out = {8'd37, 8'd110, 1'b1, 1'b0};
1479: data_out = {8'd42, 8'd110, 1'b1, 1'b0};
1480: data_out = {8'd53, 8'd110, 1'b1, 1'b0};
1481: data_out = {8'd62, 8'd110, 1'b1, 1'b0};
1482: data_out = {8'd86, 8'd110, 1'b1, 1'b0};
1483: data_out = {8'd99, 8'd110, 1'b1, 1'b0};
1484: data_out = {8'd102, 8'd110, 1'b1, 1'b0};
1485: data_out = {8'd115, 8'd110, 1'b1, 1'b0};
1486: data_out = {8'd143, 8'd110, 1'b1, 1'b0};
1487: data_out = {8'd160, 8'd110, 1'b1, 1'b0};
1488: data_out = {8'd184, 8'd110, 1'b1, 1'b0};
1489: data_out = {8'd193, 8'd110, 1'b1, 1'b0};
1490: data_out = {8'd200, 8'd110, 1'b1, 1'b0};
1491: data_out = {8'd209, 8'd110, 1'b1, 1'b0};
1492: data_out = {8'd37, 8'd111, 1'b1, 1'b0};
1493: data_out = {8'd42, 8'd111, 1'b1, 1'b0};
1494: data_out = {8'd43, 8'd111, 1'b1, 1'b0};
1495: data_out = {8'd44, 8'd111, 1'b1, 1'b0};
1496: data_out = {8'd45, 8'd111, 1'b1, 1'b0};
1497: data_out = {8'd46, 8'd111, 1'b1, 1'b0};
1498: data_out = {8'd47, 8'd111, 1'b1, 1'b0};
1499: data_out = {8'd48, 8'd111, 1'b1, 1'b0};
1500: data_out = {8'd49, 8'd111, 1'b1, 1'b0};
1501: data_out = {8'd50, 8'd111, 1'b1, 1'b0};
1502: data_out = {8'd51, 8'd111, 1'b1, 1'b0};
1503: data_out = {8'd52, 8'd111, 1'b1, 1'b0};
1504: data_out = {8'd53, 8'd111, 1'b1, 1'b0};
1505: data_out = {8'd62, 8'd111, 1'b1, 1'b0};
1506: data_out = {8'd63, 8'd111, 1'b1, 1'b0};
1507: data_out = {8'd64, 8'd111, 1'b1, 1'b0};
1508: data_out = {8'd65, 8'd111, 1'b1, 1'b0};
1509: data_out = {8'd66, 8'd111, 1'b1, 1'b0};
1510: data_out = {8'd86, 8'd111, 1'b1, 1'b0};
1511: data_out = {8'd95, 8'd111, 1'b1, 1'b0};
1512: data_out = {8'd96, 8'd111, 1'b1, 1'b0};
1513: data_out = {8'd97, 8'd111, 1'b1, 1'b0};
1514: data_out = {8'd98, 8'd111, 1'b1, 1'b0};
1515: data_out = {8'd99, 8'd111, 1'b1, 1'b0};
1516: data_out = {8'd102, 8'd111, 1'b1, 1'b0};
1517: data_out = {8'd103, 8'd111, 1'b1, 1'b0};
1518: data_out = {8'd104, 8'd111, 1'b1, 1'b0};
1519: data_out = {8'd105, 8'd111, 1'b1, 1'b0};
1520: data_out = {8'd106, 8'd111, 1'b1, 1'b0};
1521: data_out = {8'd115, 8'd111, 1'b1, 1'b0};
1522: data_out = {8'd143, 8'd111, 1'b1, 1'b0};
1523: data_out = {8'd144, 8'd111, 1'b1, 1'b0};
1524: data_out = {8'd145, 8'd111, 1'b1, 1'b0};
1525: data_out = {8'd146, 8'd111, 1'b1, 1'b0};
1526: data_out = {8'd147, 8'd111, 1'b1, 1'b0};
1527: data_out = {8'd156, 8'd111, 1'b1, 1'b0};
1528: data_out = {8'd157, 8'd111, 1'b1, 1'b0};
1529: data_out = {8'd158, 8'd111, 1'b1, 1'b0};
1530: data_out = {8'd159, 8'd111, 1'b1, 1'b0};
1531: data_out = {8'd160, 8'd111, 1'b1, 1'b0};
1532: data_out = {8'd184, 8'd111, 1'b1, 1'b0};
1533: data_out = {8'd185, 8'd111, 1'b1, 1'b0};
1534: data_out = {8'd186, 8'd111, 1'b1, 1'b0};
1535: data_out = {8'd187, 8'd111, 1'b1, 1'b0};
1536: data_out = {8'd188, 8'd111, 1'b1, 1'b0};
1537: data_out = {8'd193, 8'd111, 1'b1, 1'b0};
1538: data_out = {8'd194, 8'd111, 1'b1, 1'b0};
1539: data_out = {8'd195, 8'd111, 1'b1, 1'b0};
1540: data_out = {8'd196, 8'd111, 1'b1, 1'b0};
1541: data_out = {8'd197, 8'd111, 1'b1, 1'b0};
1542: data_out = {8'd198, 8'd111, 1'b1, 1'b0};
1543: data_out = {8'd199, 8'd111, 1'b1, 1'b0};
1544: data_out = {8'd200, 8'd111, 1'b1, 1'b0};
1545: data_out = {8'd205, 8'd111, 1'b1, 1'b0};
1546: data_out = {8'd206, 8'd111, 1'b1, 1'b0};
1547: data_out = {8'd207, 8'd111, 1'b1, 1'b0};
1548: data_out = {8'd208, 8'd111, 1'b1, 1'b0};
1549: data_out = {8'd209, 8'd111, 1'b1, 1'b0};
1550: data_out = {8'd37, 8'd112, 1'b1, 1'b0};
1551: data_out = {8'd66, 8'd112, 1'b1, 1'b0};
1552: data_out = {8'd86, 8'd112, 1'b1, 1'b0};
1553: data_out = {8'd95, 8'd112, 1'b1, 1'b0};
1554: data_out = {8'd106, 8'd112, 1'b1, 1'b0};
1555: data_out = {8'd115, 8'd112, 1'b1, 1'b0};
1556: data_out = {8'd147, 8'd112, 1'b1, 1'b0};
1557: data_out = {8'd156, 8'd112, 1'b1, 1'b0};
1558: data_out = {8'd188, 8'd112, 1'b1, 1'b0};
1559: data_out = {8'd205, 8'd112, 1'b1, 1'b0};
1560: data_out = {8'd37, 8'd113, 1'b1, 1'b0};
1561: data_out = {8'd66, 8'd113, 1'b1, 1'b0};
1562: data_out = {8'd86, 8'd113, 1'b1, 1'b0};
1563: data_out = {8'd95, 8'd113, 1'b1, 1'b0};
1564: data_out = {8'd106, 8'd113, 1'b1, 1'b0};
1565: data_out = {8'd115, 8'd113, 1'b1, 1'b0};
1566: data_out = {8'd147, 8'd113, 1'b1, 1'b0};
1567: data_out = {8'd156, 8'd113, 1'b1, 1'b0};
1568: data_out = {8'd188, 8'd113, 1'b1, 1'b0};
1569: data_out = {8'd205, 8'd113, 1'b1, 1'b0};
1570: data_out = {8'd37, 8'd114, 1'b1, 1'b0};
1571: data_out = {8'd66, 8'd114, 1'b1, 1'b0};
1572: data_out = {8'd86, 8'd114, 1'b1, 1'b0};
1573: data_out = {8'd95, 8'd114, 1'b1, 1'b0};
1574: data_out = {8'd106, 8'd114, 1'b1, 1'b0};
1575: data_out = {8'd115, 8'd114, 1'b1, 1'b0};
1576: data_out = {8'd147, 8'd114, 1'b1, 1'b0};
1577: data_out = {8'd156, 8'd114, 1'b1, 1'b0};
1578: data_out = {8'd188, 8'd114, 1'b1, 1'b0};
1579: data_out = {8'd205, 8'd114, 1'b1, 1'b0};
1580: data_out = {8'd37, 8'd115, 1'b1, 1'b0};
1581: data_out = {8'd38, 8'd115, 1'b1, 1'b0};
1582: data_out = {8'd39, 8'd115, 1'b1, 1'b0};
1583: data_out = {8'd40, 8'd115, 1'b1, 1'b0};
1584: data_out = {8'd41, 8'd115, 1'b1, 1'b0};
1585: data_out = {8'd42, 8'd115, 1'b1, 1'b0};
1586: data_out = {8'd43, 8'd115, 1'b1, 1'b0};
1587: data_out = {8'd44, 8'd115, 1'b1, 1'b0};
1588: data_out = {8'd45, 8'd115, 1'b1, 1'b0};
1589: data_out = {8'd46, 8'd115, 1'b1, 1'b0};
1590: data_out = {8'd47, 8'd115, 1'b1, 1'b0};
1591: data_out = {8'd48, 8'd115, 1'b1, 1'b0};
1592: data_out = {8'd49, 8'd115, 1'b1, 1'b0};
1593: data_out = {8'd50, 8'd115, 1'b1, 1'b0};
1594: data_out = {8'd51, 8'd115, 1'b1, 1'b0};
1595: data_out = {8'd52, 8'd115, 1'b1, 1'b0};
1596: data_out = {8'd53, 8'd115, 1'b1, 1'b0};
1597: data_out = {8'd54, 8'd115, 1'b1, 1'b0};
1598: data_out = {8'd55, 8'd115, 1'b1, 1'b0};
1599: data_out = {8'd56, 8'd115, 1'b1, 1'b0};
1600: data_out = {8'd57, 8'd115, 1'b1, 1'b0};
1601: data_out = {8'd58, 8'd115, 1'b1, 1'b0};
1602: data_out = {8'd59, 8'd115, 1'b1, 1'b0};
1603: data_out = {8'd60, 8'd115, 1'b1, 1'b0};
1604: data_out = {8'd61, 8'd115, 1'b1, 1'b0};
1605: data_out = {8'd62, 8'd115, 1'b1, 1'b0};
1606: data_out = {8'd63, 8'd115, 1'b1, 1'b0};
1607: data_out = {8'd64, 8'd115, 1'b1, 1'b0};
1608: data_out = {8'd65, 8'd115, 1'b1, 1'b0};
1609: data_out = {8'd66, 8'd115, 1'b1, 1'b0};
1610: data_out = {8'd86, 8'd115, 1'b1, 1'b0};
1611: data_out = {8'd87, 8'd115, 1'b1, 1'b0};
1612: data_out = {8'd88, 8'd115, 1'b1, 1'b0};
1613: data_out = {8'd89, 8'd115, 1'b1, 1'b0};
1614: data_out = {8'd90, 8'd115, 1'b1, 1'b0};
1615: data_out = {8'd91, 8'd115, 1'b1, 1'b0};
1616: data_out = {8'd92, 8'd115, 1'b1, 1'b0};
1617: data_out = {8'd93, 8'd115, 1'b1, 1'b0};
1618: data_out = {8'd94, 8'd115, 1'b1, 1'b0};
1619: data_out = {8'd95, 8'd115, 1'b1, 1'b0};
1620: data_out = {8'd106, 8'd115, 1'b1, 1'b0};
1621: data_out = {8'd107, 8'd115, 1'b1, 1'b0};
1622: data_out = {8'd108, 8'd115, 1'b1, 1'b0};
1623: data_out = {8'd109, 8'd115, 1'b1, 1'b0};
1624: data_out = {8'd110, 8'd115, 1'b1, 1'b0};
1625: data_out = {8'd111, 8'd115, 1'b1, 1'b0};
1626: data_out = {8'd112, 8'd115, 1'b1, 1'b0};
1627: data_out = {8'd113, 8'd115, 1'b1, 1'b0};
1628: data_out = {8'd114, 8'd115, 1'b1, 1'b0};
1629: data_out = {8'd115, 8'd115, 1'b1, 1'b0};
1630: data_out = {8'd147, 8'd115, 1'b1, 1'b0};
1631: data_out = {8'd148, 8'd115, 1'b1, 1'b0};
1632: data_out = {8'd149, 8'd115, 1'b1, 1'b0};
1633: data_out = {8'd150, 8'd115, 1'b1, 1'b0};
1634: data_out = {8'd151, 8'd115, 1'b1, 1'b0};
1635: data_out = {8'd152, 8'd115, 1'b1, 1'b0};
1636: data_out = {8'd153, 8'd115, 1'b1, 1'b0};
1637: data_out = {8'd154, 8'd115, 1'b1, 1'b0};
1638: data_out = {8'd155, 8'd115, 1'b1, 1'b0};
1639: data_out = {8'd156, 8'd115, 1'b1, 1'b0};
1640: data_out = {8'd188, 8'd115, 1'b1, 1'b0};
1641: data_out = {8'd189, 8'd115, 1'b1, 1'b0};
1642: data_out = {8'd190, 8'd115, 1'b1, 1'b0};
1643: data_out = {8'd191, 8'd115, 1'b1, 1'b0};
1644: data_out = {8'd192, 8'd115, 1'b1, 1'b0};
1645: data_out = {8'd193, 8'd115, 1'b1, 1'b0};
1646: data_out = {8'd194, 8'd115, 1'b1, 1'b0};
1647: data_out = {8'd195, 8'd115, 1'b1, 1'b0};
1648: data_out = {8'd196, 8'd115, 1'b1, 1'b0};
1649: data_out = {8'd197, 8'd115, 1'b1, 1'b0};
1650: data_out = {8'd198, 8'd115, 1'b1, 1'b0};
1651: data_out = {8'd199, 8'd115, 1'b1, 1'b0};
1652: data_out = {8'd200, 8'd115, 1'b1, 1'b0};
1653: data_out = {8'd201, 8'd115, 1'b1, 1'b0};
1654: data_out = {8'd202, 8'd115, 1'b1, 1'b0};
1655: data_out = {8'd203, 8'd115, 1'b1, 1'b0};
1656: data_out = {8'd204, 8'd115, 1'b1, 1'b0};
1657: data_out = {8'd205, 8'd115, 1'b1, 1'b0};
1658: data_out = {8'd117, 8'd140, 1'b1, 1'b0};
1659: data_out = {8'd118, 8'd140, 1'b1, 1'b0};
1660: data_out = {8'd119, 8'd140, 1'b1, 1'b0};
1661: data_out = {8'd120, 8'd140, 1'b1, 1'b0};
1662: data_out = {8'd121, 8'd140, 1'b1, 1'b0};
1663: data_out = {8'd122, 8'd140, 1'b1, 1'b0};
1664: data_out = {8'd123, 8'd140, 1'b1, 1'b0};
1665: data_out = {8'd124, 8'd140, 1'b1, 1'b0};
1666: data_out = {8'd125, 8'd140, 1'b1, 1'b0};
1667: data_out = {8'd126, 8'd140, 1'b1, 1'b0};
1668: data_out = {8'd127, 8'd140, 1'b1, 1'b0};
1669: data_out = {8'd128, 8'd140, 1'b1, 1'b0};
1670: data_out = {8'd129, 8'd140, 1'b1, 1'b0};
1671: data_out = {8'd130, 8'd140, 1'b1, 1'b0};
1672: data_out = {8'd131, 8'd140, 1'b1, 1'b0};
1673: data_out = {8'd132, 8'd140, 1'b1, 1'b0};
1674: data_out = {8'd133, 8'd140, 1'b1, 1'b0};
1675: data_out = {8'd134, 8'd140, 1'b1, 1'b0};
1676: data_out = {8'd135, 8'd140, 1'b1, 1'b0};
1677: data_out = {8'd136, 8'd140, 1'b1, 1'b0};
1678: data_out = {8'd137, 8'd140, 1'b1, 1'b0};
1679: data_out = {8'd113, 8'd141, 1'b1, 1'b0};
1680: data_out = {8'd114, 8'd141, 1'b1, 1'b0};
1681: data_out = {8'd115, 8'd141, 1'b1, 1'b0};
1682: data_out = {8'd116, 8'd141, 1'b1, 1'b0};
1683: data_out = {8'd117, 8'd141, 1'b1, 1'b0};
1684: data_out = {8'd137, 8'd141, 1'b1, 1'b0};
1685: data_out = {8'd138, 8'd141, 1'b1, 1'b0};
1686: data_out = {8'd139, 8'd141, 1'b1, 1'b0};
1687: data_out = {8'd140, 8'd141, 1'b1, 1'b0};
1688: data_out = {8'd141, 8'd141, 1'b1, 1'b0};
1689: data_out = {8'd110, 8'd142, 1'b1, 1'b0};
1690: data_out = {8'd111, 8'd142, 1'b1, 1'b0};
1691: data_out = {8'd112, 8'd142, 1'b1, 1'b0};
1692: data_out = {8'd113, 8'd142, 1'b1, 1'b0};
1693: data_out = {8'd141, 8'd142, 1'b1, 1'b0};
1694: data_out = {8'd142, 8'd142, 1'b1, 1'b0};
1695: data_out = {8'd143, 8'd142, 1'b1, 1'b0};
1696: data_out = {8'd144, 8'd142, 1'b1, 1'b0};
1697: data_out = {8'd108, 8'd143, 1'b1, 1'b0};
1698: data_out = {8'd109, 8'd143, 1'b1, 1'b0};
1699: data_out = {8'd110, 8'd143, 1'b1, 1'b0};
1700: data_out = {8'd144, 8'd143, 1'b1, 1'b0};
1701: data_out = {8'd145, 8'd143, 1'b1, 1'b0};
1702: data_out = {8'd146, 8'd143, 1'b1, 1'b0};
1703: data_out = {8'd105, 8'd144, 1'b1, 1'b0};
1704: data_out = {8'd106, 8'd144, 1'b1, 1'b0};
1705: data_out = {8'd107, 8'd144, 1'b1, 1'b0};
1706: data_out = {8'd108, 8'd144, 1'b1, 1'b0};
1707: data_out = {8'd146, 8'd144, 1'b1, 1'b0};
1708: data_out = {8'd147, 8'd144, 1'b1, 1'b0};
1709: data_out = {8'd148, 8'd144, 1'b1, 1'b0};
1710: data_out = {8'd149, 8'd144, 1'b1, 1'b0};
1711: data_out = {8'd103, 8'd145, 1'b1, 1'b0};
1712: data_out = {8'd104, 8'd145, 1'b1, 1'b0};
1713: data_out = {8'd105, 8'd145, 1'b1, 1'b0};
1714: data_out = {8'd149, 8'd145, 1'b1, 1'b0};
1715: data_out = {8'd150, 8'd145, 1'b1, 1'b0};
1716: data_out = {8'd151, 8'd145, 1'b1, 1'b0};
1717: data_out = {8'd102, 8'd146, 1'b1, 1'b0};
1718: data_out = {8'd103, 8'd146, 1'b1, 1'b0};
1719: data_out = {8'd151, 8'd146, 1'b1, 1'b0};
1720: data_out = {8'd152, 8'd146, 1'b1, 1'b0};
1721: data_out = {8'd102, 8'd147, 1'b1, 1'b0};
1722: data_out = {8'd152, 8'd147, 1'b1, 1'b0};
1723: data_out = {8'd102, 8'd148, 1'b1, 1'b0};
1724: data_out = {8'd103, 8'd148, 1'b1, 1'b0};
1725: data_out = {8'd151, 8'd148, 1'b1, 1'b0};
1726: data_out = {8'd152, 8'd148, 1'b1, 1'b0};
1727: data_out = {8'd103, 8'd149, 1'b1, 1'b0};
1728: data_out = {8'd104, 8'd149, 1'b1, 1'b0};
1729: data_out = {8'd150, 8'd149, 1'b1, 1'b0};
1730: data_out = {8'd151, 8'd149, 1'b1, 1'b0};
1731: data_out = {8'd104, 8'd150, 1'b1, 1'b0};
1732: data_out = {8'd150, 8'd150, 1'b1, 1'b0};
1733: data_out = {8'd104, 8'd151, 1'b1, 1'b0};
1734: data_out = {8'd105, 8'd151, 1'b1, 1'b0};
1735: data_out = {8'd149, 8'd151, 1'b1, 1'b0};
1736: data_out = {8'd150, 8'd151, 1'b1, 1'b0};
1737: data_out = {8'd105, 8'd152, 1'b1, 1'b0};
1738: data_out = {8'd149, 8'd152, 1'b1, 1'b0};
1739: data_out = {8'd105, 8'd153, 1'b1, 1'b0};
1740: data_out = {8'd106, 8'd153, 1'b1, 1'b0};
1741: data_out = {8'd148, 8'd153, 1'b1, 1'b0};
1742: data_out = {8'd149, 8'd153, 1'b1, 1'b0};
1743: data_out = {8'd106, 8'd154, 1'b1, 1'b0};
1744: data_out = {8'd148, 8'd154, 1'b1, 1'b0};
1745: data_out = {8'd106, 8'd155, 1'b1, 1'b0};
1746: data_out = {8'd107, 8'd155, 1'b1, 1'b0};
1747: data_out = {8'd147, 8'd155, 1'b1, 1'b0};
1748: data_out = {8'd148, 8'd155, 1'b1, 1'b0};
1749: data_out = {8'd107, 8'd156, 1'b1, 1'b0};
1750: data_out = {8'd108, 8'd156, 1'b1, 1'b0};
1751: data_out = {8'd146, 8'd156, 1'b1, 1'b0};
1752: data_out = {8'd147, 8'd156, 1'b1, 1'b0};
1753: data_out = {8'd108, 8'd157, 1'b1, 1'b0};
1754: data_out = {8'd146, 8'd157, 1'b1, 1'b0};
1755: data_out = {8'd108, 8'd158, 1'b1, 1'b0};
1756: data_out = {8'd109, 8'd158, 1'b1, 1'b0};
1757: data_out = {8'd145, 8'd158, 1'b1, 1'b0};
1758: data_out = {8'd146, 8'd158, 1'b1, 1'b0};
1759: data_out = {8'd109, 8'd159, 1'b1, 1'b0};
1760: data_out = {8'd145, 8'd159, 1'b1, 1'b0};
1761: data_out = {8'd109, 8'd160, 1'b1, 1'b0};
1762: data_out = {8'd110, 8'd160, 1'b1, 1'b0};
1763: data_out = {8'd144, 8'd160, 1'b1, 1'b0};
1764: data_out = {8'd145, 8'd160, 1'b1, 1'b0};
1765: data_out = {8'd110, 8'd161, 1'b1, 1'b0};
1766: data_out = {8'd144, 8'd161, 1'b1, 1'b0};
1767: data_out = {8'd110, 8'd162, 1'b1, 1'b0};
1768: data_out = {8'd111, 8'd162, 1'b1, 1'b0};
1769: data_out = {8'd143, 8'd162, 1'b1, 1'b0};
1770: data_out = {8'd144, 8'd162, 1'b1, 1'b0};
1771: data_out = {8'd111, 8'd163, 1'b1, 1'b0};
1772: data_out = {8'd112, 8'd163, 1'b1, 1'b0};
1773: data_out = {8'd142, 8'd163, 1'b1, 1'b0};
1774: data_out = {8'd143, 8'd163, 1'b1, 1'b0};
1775: data_out = {8'd112, 8'd164, 1'b1, 1'b0};
1776: data_out = {8'd142, 8'd164, 1'b1, 1'b0};
1777: data_out = {8'd112, 8'd165, 1'b1, 1'b0};
1778: data_out = {8'd113, 8'd165, 1'b1, 1'b0};
1779: data_out = {8'd141, 8'd165, 1'b1, 1'b0};
1780: data_out = {8'd142, 8'd165, 1'b1, 1'b0};
1781: data_out = {8'd113, 8'd166, 1'b1, 1'b0};
1782: data_out = {8'd141, 8'd166, 1'b1, 1'b0};
1783: data_out = {8'd113, 8'd167, 1'b1, 1'b0};
1784: data_out = {8'd114, 8'd167, 1'b1, 1'b0};
1785: data_out = {8'd140, 8'd167, 1'b1, 1'b0};
1786: data_out = {8'd141, 8'd167, 1'b1, 1'b0};
1787: data_out = {8'd114, 8'd168, 1'b1, 1'b0};
1788: data_out = {8'd115, 8'd168, 1'b1, 1'b0};
1789: data_out = {8'd139, 8'd168, 1'b1, 1'b0};
1790: data_out = {8'd140, 8'd168, 1'b1, 1'b0};
1791: data_out = {8'd115, 8'd169, 1'b1, 1'b0};
1792: data_out = {8'd139, 8'd169, 1'b1, 1'b0};
1793: data_out = {8'd115, 8'd170, 1'b1, 1'b0};
1794: data_out = {8'd116, 8'd170, 1'b1, 1'b0};
1795: data_out = {8'd138, 8'd170, 1'b1, 1'b0};
1796: data_out = {8'd139, 8'd170, 1'b1, 1'b0};
1797: data_out = {8'd116, 8'd171, 1'b1, 1'b0};
1798: data_out = {8'd138, 8'd171, 1'b1, 1'b0};
1799: data_out = {8'd116, 8'd172, 1'b1, 1'b0};
1800: data_out = {8'd117, 8'd172, 1'b1, 1'b0};
1801: data_out = {8'd137, 8'd172, 1'b1, 1'b0};
1802: data_out = {8'd138, 8'd172, 1'b1, 1'b0};
1803: data_out = {8'd117, 8'd173, 1'b1, 1'b0};
1804: data_out = {8'd137, 8'd173, 1'b1, 1'b0};
1805: data_out = {8'd117, 8'd174, 1'b1, 1'b0};
1806: data_out = {8'd118, 8'd174, 1'b1, 1'b0};
1807: data_out = {8'd136, 8'd174, 1'b1, 1'b0};
1808: data_out = {8'd137, 8'd174, 1'b1, 1'b0};
1809: data_out = {8'd118, 8'd175, 1'b1, 1'b0};
1810: data_out = {8'd119, 8'd175, 1'b1, 1'b0};
1811: data_out = {8'd124, 8'd175, 1'b1, 1'b0};
1812: data_out = {8'd125, 8'd175, 1'b1, 1'b0};
1813: data_out = {8'd126, 8'd175, 1'b1, 1'b0};
1814: data_out = {8'd127, 8'd175, 1'b1, 1'b0};
1815: data_out = {8'd128, 8'd175, 1'b1, 1'b0};
1816: data_out = {8'd129, 8'd175, 1'b1, 1'b0};
1817: data_out = {8'd130, 8'd175, 1'b1, 1'b0};
1818: data_out = {8'd135, 8'd175, 1'b1, 1'b0};
1819: data_out = {8'd136, 8'd175, 1'b1, 1'b0};
1820: data_out = {8'd119, 8'd176, 1'b1, 1'b0};
1821: data_out = {8'd120, 8'd176, 1'b1, 1'b0};
1822: data_out = {8'd121, 8'd176, 1'b1, 1'b0};
1823: data_out = {8'd122, 8'd176, 1'b1, 1'b0};
1824: data_out = {8'd123, 8'd176, 1'b1, 1'b0};
1825: data_out = {8'd124, 8'd176, 1'b1, 1'b0};
1826: data_out = {8'd130, 8'd176, 1'b1, 1'b0};
1827: data_out = {8'd131, 8'd176, 1'b1, 1'b0};
1828: data_out = {8'd132, 8'd176, 1'b1, 1'b0};
1829: data_out = {8'd133, 8'd176, 1'b1, 1'b0};
1830: data_out = {8'd134, 8'd176, 1'b1, 1'b0};
1831: data_out = {8'd135, 8'd176, 1'b1, 1'b0};
1832: data_out = {8'd119, 8'd177, 1'b1, 1'b0};
1833: data_out = {8'd120, 8'd177, 1'b1, 1'b0};
1834: data_out = {8'd134, 8'd177, 1'b1, 1'b0};
1835: data_out = {8'd135, 8'd177, 1'b1, 1'b0};
1836: data_out = {8'd124, 8'd181, 1'b1, 1'b0};
1837: data_out = {8'd125, 8'd181, 1'b1, 1'b0};
1838: data_out = {8'd126, 8'd181, 1'b1, 1'b0};
1839: data_out = {8'd127, 8'd181, 1'b1, 1'b0};
1840: data_out = {8'd128, 8'd181, 1'b1, 1'b0};
1841: data_out = {8'd129, 8'd181, 1'b1, 1'b0};
1842: data_out = {8'd130, 8'd181, 1'b1, 1'b0};
1843: data_out = {8'd122, 8'd182, 1'b1, 1'b0};
1844: data_out = {8'd123, 8'd182, 1'b1, 1'b0};
1845: data_out = {8'd124, 8'd182, 1'b1, 1'b0};
1846: data_out = {8'd130, 8'd182, 1'b1, 1'b0};
1847: data_out = {8'd131, 8'd182, 1'b1, 1'b0};
1848: data_out = {8'd132, 8'd182, 1'b1, 1'b0};
1849: data_out = {8'd121, 8'd183, 1'b1, 1'b0};
1850: data_out = {8'd122, 8'd183, 1'b1, 1'b0};
1851: data_out = {8'd132, 8'd183, 1'b1, 1'b0};
1852: data_out = {8'd133, 8'd183, 1'b1, 1'b0};
1853: data_out = {8'd120, 8'd184, 1'b1, 1'b0};
1854: data_out = {8'd121, 8'd184, 1'b1, 1'b0};
1855: data_out = {8'd133, 8'd184, 1'b1, 1'b0};
1856: data_out = {8'd134, 8'd184, 1'b1, 1'b0};
1857: data_out = {8'd119, 8'd185, 1'b1, 1'b0};
1858: data_out = {8'd120, 8'd185, 1'b1, 1'b0};
1859: data_out = {8'd134, 8'd185, 1'b1, 1'b0};
1860: data_out = {8'd135, 8'd185, 1'b1, 1'b0};
1861: data_out = {8'd118, 8'd186, 1'b1, 1'b0};
1862: data_out = {8'd119, 8'd186, 1'b1, 1'b0};
1863: data_out = {8'd135, 8'd186, 1'b1, 1'b0};
1864: data_out = {8'd136, 8'd186, 1'b1, 1'b0};
1865: data_out = {8'd118, 8'd187, 1'b1, 1'b0};
1866: data_out = {8'd136, 8'd187, 1'b1, 1'b0};
1867: data_out = {8'd117, 8'd188, 1'b1, 1'b0};
1868: data_out = {8'd118, 8'd188, 1'b1, 1'b0};
1869: data_out = {8'd136, 8'd188, 1'b1, 1'b0};
1870: data_out = {8'd137, 8'd188, 1'b1, 1'b0};
1871: data_out = {8'd117, 8'd189, 1'b1, 1'b0};
1872: data_out = {8'd137, 8'd189, 1'b1, 1'b0};
1873: data_out = {8'd117, 8'd190, 1'b1, 1'b0};
1874: data_out = {8'd137, 8'd190, 1'b1, 1'b0};
1875: data_out = {8'd76, 8'd191, 1'b1, 1'b0};
1876: data_out = {8'd77, 8'd191, 1'b1, 1'b0};
1877: data_out = {8'd78, 8'd191, 1'b1, 1'b0};
1878: data_out = {8'd79, 8'd191, 1'b1, 1'b0};
1879: data_out = {8'd80, 8'd191, 1'b1, 1'b0};
1880: data_out = {8'd81, 8'd191, 1'b1, 1'b0};
1881: data_out = {8'd82, 8'd191, 1'b1, 1'b0};
1882: data_out = {8'd83, 8'd191, 1'b1, 1'b0};
1883: data_out = {8'd84, 8'd191, 1'b1, 1'b0};
1884: data_out = {8'd85, 8'd191, 1'b1, 1'b0};
1885: data_out = {8'd86, 8'd191, 1'b1, 1'b0};
1886: data_out = {8'd87, 8'd191, 1'b1, 1'b0};
1887: data_out = {8'd88, 8'd191, 1'b1, 1'b0};
1888: data_out = {8'd89, 8'd191, 1'b1, 1'b0};
1889: data_out = {8'd90, 8'd191, 1'b1, 1'b0};
1890: data_out = {8'd91, 8'd191, 1'b1, 1'b0};
1891: data_out = {8'd92, 8'd191, 1'b1, 1'b0};
1892: data_out = {8'd93, 8'd191, 1'b1, 1'b0};
1893: data_out = {8'd94, 8'd191, 1'b1, 1'b0};
1894: data_out = {8'd95, 8'd191, 1'b1, 1'b0};
1895: data_out = {8'd96, 8'd191, 1'b1, 1'b0};
1896: data_out = {8'd97, 8'd191, 1'b1, 1'b0};
1897: data_out = {8'd98, 8'd191, 1'b1, 1'b0};
1898: data_out = {8'd99, 8'd191, 1'b1, 1'b0};
1899: data_out = {8'd100, 8'd191, 1'b1, 1'b0};
1900: data_out = {8'd101, 8'd191, 1'b1, 1'b0};
1901: data_out = {8'd102, 8'd191, 1'b1, 1'b0};
1902: data_out = {8'd103, 8'd191, 1'b1, 1'b0};
1903: data_out = {8'd104, 8'd191, 1'b1, 1'b0};
1904: data_out = {8'd105, 8'd191, 1'b1, 1'b0};
1905: data_out = {8'd106, 8'd191, 1'b1, 1'b0};
1906: data_out = {8'd107, 8'd191, 1'b1, 1'b0};
1907: data_out = {8'd108, 8'd191, 1'b1, 1'b0};
1908: data_out = {8'd109, 8'd191, 1'b1, 1'b0};
1909: data_out = {8'd110, 8'd191, 1'b1, 1'b0};
1910: data_out = {8'd111, 8'd191, 1'b1, 1'b0};
1911: data_out = {8'd117, 8'd191, 1'b1, 1'b0};
1912: data_out = {8'd137, 8'd191, 1'b1, 1'b0};
1913: data_out = {8'd143, 8'd191, 1'b1, 1'b0};
1914: data_out = {8'd144, 8'd191, 1'b1, 1'b0};
1915: data_out = {8'd145, 8'd191, 1'b1, 1'b0};
1916: data_out = {8'd146, 8'd191, 1'b1, 1'b0};
1917: data_out = {8'd147, 8'd191, 1'b1, 1'b0};
1918: data_out = {8'd148, 8'd191, 1'b1, 1'b0};
1919: data_out = {8'd149, 8'd191, 1'b1, 1'b0};
1920: data_out = {8'd150, 8'd191, 1'b1, 1'b0};
1921: data_out = {8'd151, 8'd191, 1'b1, 1'b0};
1922: data_out = {8'd152, 8'd191, 1'b1, 1'b0};
1923: data_out = {8'd153, 8'd191, 1'b1, 1'b0};
1924: data_out = {8'd154, 8'd191, 1'b1, 1'b0};
1925: data_out = {8'd155, 8'd191, 1'b1, 1'b0};
1926: data_out = {8'd156, 8'd191, 1'b1, 1'b0};
1927: data_out = {8'd157, 8'd191, 1'b1, 1'b0};
1928: data_out = {8'd158, 8'd191, 1'b1, 1'b0};
1929: data_out = {8'd159, 8'd191, 1'b1, 1'b0};
1930: data_out = {8'd160, 8'd191, 1'b1, 1'b0};
1931: data_out = {8'd161, 8'd191, 1'b1, 1'b0};
1932: data_out = {8'd162, 8'd191, 1'b1, 1'b0};
1933: data_out = {8'd163, 8'd191, 1'b1, 1'b0};
1934: data_out = {8'd164, 8'd191, 1'b1, 1'b0};
1935: data_out = {8'd165, 8'd191, 1'b1, 1'b0};
1936: data_out = {8'd166, 8'd191, 1'b1, 1'b0};
1937: data_out = {8'd167, 8'd191, 1'b1, 1'b0};
1938: data_out = {8'd168, 8'd191, 1'b1, 1'b0};
1939: data_out = {8'd169, 8'd191, 1'b1, 1'b0};
1940: data_out = {8'd170, 8'd191, 1'b1, 1'b0};
1941: data_out = {8'd171, 8'd191, 1'b1, 1'b0};
1942: data_out = {8'd172, 8'd191, 1'b1, 1'b0};
1943: data_out = {8'd173, 8'd191, 1'b1, 1'b0};
1944: data_out = {8'd174, 8'd191, 1'b1, 1'b0};
1945: data_out = {8'd175, 8'd191, 1'b1, 1'b0};
1946: data_out = {8'd176, 8'd191, 1'b1, 1'b0};
1947: data_out = {8'd177, 8'd191, 1'b1, 1'b0};
1948: data_out = {8'd178, 8'd191, 1'b1, 1'b0};
1949: data_out = {8'd76, 8'd192, 1'b1, 1'b0};
1950: data_out = {8'd111, 8'd192, 1'b1, 1'b0};
1951: data_out = {8'd117, 8'd192, 1'b1, 1'b0};
1952: data_out = {8'd137, 8'd192, 1'b1, 1'b0};
1953: data_out = {8'd143, 8'd192, 1'b1, 1'b0};
1954: data_out = {8'd178, 8'd192, 1'b1, 1'b0};
1955: data_out = {8'd179, 8'd192, 1'b1, 1'b0};
1956: data_out = {8'd76, 8'd193, 1'b1, 1'b0};
1957: data_out = {8'd111, 8'd193, 1'b1, 1'b0};
1958: data_out = {8'd117, 8'd193, 1'b1, 1'b0};
1959: data_out = {8'd137, 8'd193, 1'b1, 1'b0};
1960: data_out = {8'd143, 8'd193, 1'b1, 1'b0};
1961: data_out = {8'd178, 8'd193, 1'b1, 1'b0};
1962: data_out = {8'd76, 8'd194, 1'b1, 1'b0};
1963: data_out = {8'd111, 8'd194, 1'b1, 1'b0};
1964: data_out = {8'd112, 8'd194, 1'b1, 1'b0};
1965: data_out = {8'd117, 8'd194, 1'b1, 1'b0};
1966: data_out = {8'd118, 8'd194, 1'b1, 1'b0};
1967: data_out = {8'd136, 8'd194, 1'b1, 1'b0};
1968: data_out = {8'd137, 8'd194, 1'b1, 1'b0};
1969: data_out = {8'd142, 8'd194, 1'b1, 1'b0};
1970: data_out = {8'd143, 8'd194, 1'b1, 1'b0};
1971: data_out = {8'd178, 8'd194, 1'b1, 1'b0};
1972: data_out = {8'd76, 8'd195, 1'b1, 1'b0};
1973: data_out = {8'd112, 8'd195, 1'b1, 1'b0};
1974: data_out = {8'd118, 8'd195, 1'b1, 1'b0};
1975: data_out = {8'd136, 8'd195, 1'b1, 1'b0};
1976: data_out = {8'd142, 8'd195, 1'b1, 1'b0};
1977: data_out = {8'd178, 8'd195, 1'b1, 1'b0};
1978: data_out = {8'd76, 8'd196, 1'b1, 1'b0};
1979: data_out = {8'd112, 8'd196, 1'b1, 1'b0};
1980: data_out = {8'd118, 8'd196, 1'b1, 1'b0};
1981: data_out = {8'd119, 8'd196, 1'b1, 1'b0};
1982: data_out = {8'd135, 8'd196, 1'b1, 1'b0};
1983: data_out = {8'd136, 8'd196, 1'b1, 1'b0};
1984: data_out = {8'd142, 8'd196, 1'b1, 1'b0};
1985: data_out = {8'd178, 8'd196, 1'b1, 1'b0};
1986: data_out = {8'd76, 8'd197, 1'b1, 1'b0};
1987: data_out = {8'd112, 8'd197, 1'b1, 1'b0};
1988: data_out = {8'd119, 8'd197, 1'b1, 1'b0};
1989: data_out = {8'd120, 8'd197, 1'b1, 1'b0};
1990: data_out = {8'd134, 8'd197, 1'b1, 1'b0};
1991: data_out = {8'd135, 8'd197, 1'b1, 1'b0};
1992: data_out = {8'd142, 8'd197, 1'b1, 1'b0};
1993: data_out = {8'd178, 8'd197, 1'b1, 1'b0};
1994: data_out = {8'd76, 8'd198, 1'b1, 1'b0};
1995: data_out = {8'd112, 8'd198, 1'b1, 1'b0};
1996: data_out = {8'd113, 8'd198, 1'b1, 1'b0};
1997: data_out = {8'd120, 8'd198, 1'b1, 1'b0};
1998: data_out = {8'd121, 8'd198, 1'b1, 1'b0};
1999: data_out = {8'd133, 8'd198, 1'b1, 1'b0};
2000: data_out = {8'd134, 8'd198, 1'b1, 1'b0};
2001: data_out = {8'd141, 8'd198, 1'b1, 1'b0};
2002: data_out = {8'd142, 8'd198, 1'b1, 1'b0};
2003: data_out = {8'd178, 8'd198, 1'b1, 1'b0};
2004: data_out = {8'd76, 8'd199, 1'b1, 1'b0};
2005: data_out = {8'd113, 8'd199, 1'b1, 1'b0};
2006: data_out = {8'd121, 8'd199, 1'b1, 1'b0};
2007: data_out = {8'd122, 8'd199, 1'b1, 1'b0};
2008: data_out = {8'd132, 8'd199, 1'b1, 1'b0};
2009: data_out = {8'd133, 8'd199, 1'b1, 1'b0};
2010: data_out = {8'd141, 8'd199, 1'b1, 1'b0};
2011: data_out = {8'd178, 8'd199, 1'b1, 1'b0};
2012: data_out = {8'd76, 8'd200, 1'b1, 1'b0};
2013: data_out = {8'd113, 8'd200, 1'b1, 1'b0};
2014: data_out = {8'd114, 8'd200, 1'b1, 1'b0};
2015: data_out = {8'd122, 8'd200, 1'b1, 1'b0};
2016: data_out = {8'd123, 8'd200, 1'b1, 1'b0};
2017: data_out = {8'd124, 8'd200, 1'b1, 1'b0};
2018: data_out = {8'd130, 8'd200, 1'b1, 1'b0};
2019: data_out = {8'd131, 8'd200, 1'b1, 1'b0};
2020: data_out = {8'd132, 8'd200, 1'b1, 1'b0};
2021: data_out = {8'd140, 8'd200, 1'b1, 1'b0};
2022: data_out = {8'd141, 8'd200, 1'b1, 1'b0};
2023: data_out = {8'd178, 8'd200, 1'b1, 1'b0};
2024: data_out = {8'd76, 8'd201, 1'b1, 1'b0};
2025: data_out = {8'd77, 8'd201, 1'b1, 1'b0};
2026: data_out = {8'd114, 8'd201, 1'b1, 1'b0};
2027: data_out = {8'd115, 8'd201, 1'b1, 1'b0};
2028: data_out = {8'd124, 8'd201, 1'b1, 1'b0};
2029: data_out = {8'd125, 8'd201, 1'b1, 1'b0};
2030: data_out = {8'd126, 8'd201, 1'b1, 1'b0};
2031: data_out = {8'd127, 8'd201, 1'b1, 1'b0};
2032: data_out = {8'd128, 8'd201, 1'b1, 1'b0};
2033: data_out = {8'd129, 8'd201, 1'b1, 1'b0};
2034: data_out = {8'd130, 8'd201, 1'b1, 1'b0};
2035: data_out = {8'd139, 8'd201, 1'b1, 1'b0};
2036: data_out = {8'd140, 8'd201, 1'b1, 1'b0};
2037: data_out = {8'd177, 8'd201, 1'b1, 1'b0};
2038: data_out = {8'd178, 8'd201, 1'b1, 1'b0};
2039: data_out = {8'd77, 8'd202, 1'b1, 1'b0};
2040: data_out = {8'd115, 8'd202, 1'b1, 1'b0};
2041: data_out = {8'd116, 8'd202, 1'b1, 1'b0};
2042: data_out = {8'd138, 8'd202, 1'b1, 1'b0};
2043: data_out = {8'd139, 8'd202, 1'b1, 1'b0};
2044: data_out = {8'd177, 8'd202, 1'b1, 1'b0};
2045: data_out = {8'd77, 8'd203, 1'b1, 1'b0};
2046: data_out = {8'd116, 8'd203, 1'b1, 1'b0};
2047: data_out = {8'd117, 8'd203, 1'b1, 1'b0};
2048: data_out = {8'd137, 8'd203, 1'b1, 1'b0};
2049: data_out = {8'd138, 8'd203, 1'b1, 1'b0};
2050: data_out = {8'd177, 8'd203, 1'b1, 1'b0};
2051: data_out = {8'd77, 8'd204, 1'b1, 1'b0};
2052: data_out = {8'd117, 8'd204, 1'b1, 1'b0};
2053: data_out = {8'd118, 8'd204, 1'b1, 1'b0};
2054: data_out = {8'd136, 8'd204, 1'b1, 1'b0};
2055: data_out = {8'd137, 8'd204, 1'b1, 1'b0};
2056: data_out = {8'd177, 8'd204, 1'b1, 1'b0};
2057: data_out = {8'd77, 8'd205, 1'b1, 1'b0};
2058: data_out = {8'd78, 8'd205, 1'b1, 1'b0};
2059: data_out = {8'd118, 8'd205, 1'b1, 1'b0};
2060: data_out = {8'd119, 8'd205, 1'b1, 1'b0};
2061: data_out = {8'd135, 8'd205, 1'b1, 1'b0};
2062: data_out = {8'd136, 8'd205, 1'b1, 1'b0};
2063: data_out = {8'd176, 8'd205, 1'b1, 1'b0};
2064: data_out = {8'd177, 8'd205, 1'b1, 1'b0};
2065: data_out = {8'd78, 8'd206, 1'b1, 1'b0};
2066: data_out = {8'd118, 8'd206, 1'b1, 1'b0};
2067: data_out = {8'd136, 8'd206, 1'b1, 1'b0};
2068: data_out = {8'd176, 8'd206, 1'b1, 1'b0};
2069: data_out = {8'd78, 8'd207, 1'b1, 1'b0};
2070: data_out = {8'd117, 8'd207, 1'b1, 1'b0};
2071: data_out = {8'd118, 8'd207, 1'b1, 1'b0};
2072: data_out = {8'd136, 8'd207, 1'b1, 1'b0};
2073: data_out = {8'd137, 8'd207, 1'b1, 1'b0};
2074: data_out = {8'd176, 8'd207, 1'b1, 1'b0};
2075: data_out = {8'd78, 8'd208, 1'b1, 1'b0};
2076: data_out = {8'd79, 8'd208, 1'b1, 1'b0};
2077: data_out = {8'd116, 8'd208, 1'b1, 1'b0};
2078: data_out = {8'd117, 8'd208, 1'b1, 1'b0};
2079: data_out = {8'd137, 8'd208, 1'b1, 1'b0};
2080: data_out = {8'd138, 8'd208, 1'b1, 1'b0};
2081: data_out = {8'd175, 8'd208, 1'b1, 1'b0};
2082: data_out = {8'd176, 8'd208, 1'b1, 1'b0};
2083: data_out = {8'd79, 8'd209, 1'b1, 1'b0};
2084: data_out = {8'd116, 8'd209, 1'b1, 1'b0};
2085: data_out = {8'd138, 8'd209, 1'b1, 1'b0};
2086: data_out = {8'd175, 8'd209, 1'b1, 1'b0};
2087: data_out = {8'd79, 8'd210, 1'b1, 1'b0};
2088: data_out = {8'd115, 8'd210, 1'b1, 1'b0};
2089: data_out = {8'd116, 8'd210, 1'b1, 1'b0};
2090: data_out = {8'd138, 8'd210, 1'b1, 1'b0};
2091: data_out = {8'd139, 8'd210, 1'b1, 1'b0};
2092: data_out = {8'd175, 8'd210, 1'b1, 1'b0};
2093: data_out = {8'd79, 8'd211, 1'b1, 1'b0};
2094: data_out = {8'd80, 8'd211, 1'b1, 1'b0};
2095: data_out = {8'd115, 8'd211, 1'b1, 1'b0};
2096: data_out = {8'd139, 8'd211, 1'b1, 1'b0};
2097: data_out = {8'd174, 8'd211, 1'b1, 1'b0};
2098: data_out = {8'd175, 8'd211, 1'b1, 1'b0};
2099: data_out = {8'd80, 8'd212, 1'b1, 1'b0};
2100: data_out = {8'd114, 8'd212, 1'b1, 1'b0};
2101: data_out = {8'd115, 8'd212, 1'b1, 1'b0};
2102: data_out = {8'd139, 8'd212, 1'b1, 1'b0};
2103: data_out = {8'd140, 8'd212, 1'b1, 1'b0};
2104: data_out = {8'd174, 8'd212, 1'b1, 1'b0};
2105: data_out = {8'd80, 8'd213, 1'b1, 1'b0};
2106: data_out = {8'd81, 8'd213, 1'b1, 1'b0};
2107: data_out = {8'd113, 8'd213, 1'b1, 1'b0};
2108: data_out = {8'd114, 8'd213, 1'b1, 1'b0};
2109: data_out = {8'd140, 8'd213, 1'b1, 1'b0};
2110: data_out = {8'd141, 8'd213, 1'b1, 1'b0};
2111: data_out = {8'd173, 8'd213, 1'b1, 1'b0};
2112: data_out = {8'd174, 8'd213, 1'b1, 1'b0};
2113: data_out = {8'd81, 8'd214, 1'b1, 1'b0};
2114: data_out = {8'd113, 8'd214, 1'b1, 1'b0};
2115: data_out = {8'd141, 8'd214, 1'b1, 1'b0};
2116: data_out = {8'd173, 8'd214, 1'b1, 1'b0};
2117: data_out = {8'd81, 8'd215, 1'b1, 1'b0};
2118: data_out = {8'd82, 8'd215, 1'b1, 1'b0};
2119: data_out = {8'd112, 8'd215, 1'b1, 1'b0};
2120: data_out = {8'd113, 8'd215, 1'b1, 1'b0};
2121: data_out = {8'd141, 8'd215, 1'b1, 1'b0};
2122: data_out = {8'd142, 8'd215, 1'b1, 1'b0};
2123: data_out = {8'd172, 8'd215, 1'b1, 1'b0};
2124: data_out = {8'd173, 8'd215, 1'b1, 1'b0};
2125: data_out = {8'd82, 8'd216, 1'b1, 1'b0};
2126: data_out = {8'd112, 8'd216, 1'b1, 1'b0};
2127: data_out = {8'd142, 8'd216, 1'b1, 1'b0};
2128: data_out = {8'd172, 8'd216, 1'b1, 1'b0};
2129: data_out = {8'd82, 8'd217, 1'b1, 1'b0};
2130: data_out = {8'd83, 8'd217, 1'b1, 1'b0};
2131: data_out = {8'd111, 8'd217, 1'b1, 1'b0};
2132: data_out = {8'd112, 8'd217, 1'b1, 1'b0};
2133: data_out = {8'd142, 8'd217, 1'b1, 1'b0};
2134: data_out = {8'd143, 8'd217, 1'b1, 1'b0};
2135: data_out = {8'd171, 8'd217, 1'b1, 1'b0};
2136: data_out = {8'd172, 8'd217, 1'b1, 1'b0};
2137: data_out = {8'd83, 8'd218, 1'b1, 1'b0};
2138: data_out = {8'd84, 8'd218, 1'b1, 1'b0};
2139: data_out = {8'd111, 8'd218, 1'b1, 1'b0};
2140: data_out = {8'd143, 8'd218, 1'b1, 1'b0};
2141: data_out = {8'd170, 8'd218, 1'b1, 1'b0};
2142: data_out = {8'd171, 8'd218, 1'b1, 1'b0};
2143: data_out = {8'd84, 8'd219, 1'b1, 1'b0};
2144: data_out = {8'd110, 8'd219, 1'b1, 1'b0};
2145: data_out = {8'd111, 8'd219, 1'b1, 1'b0};
2146: data_out = {8'd143, 8'd219, 1'b1, 1'b0};
2147: data_out = {8'd144, 8'd219, 1'b1, 1'b0};
2148: data_out = {8'd170, 8'd219, 1'b1, 1'b0};
2149: data_out = {8'd84, 8'd220, 1'b1, 1'b0};
2150: data_out = {8'd85, 8'd220, 1'b1, 1'b0};
2151: data_out = {8'd109, 8'd220, 1'b1, 1'b0};
2152: data_out = {8'd110, 8'd220, 1'b1, 1'b0};
2153: data_out = {8'd144, 8'd220, 1'b1, 1'b0};
2154: data_out = {8'd145, 8'd220, 1'b1, 1'b0};
2155: data_out = {8'd169, 8'd220, 1'b1, 1'b0};
2156: data_out = {8'd170, 8'd220, 1'b1, 1'b0};
2157: data_out = {8'd85, 8'd221, 1'b1, 1'b0};
2158: data_out = {8'd86, 8'd221, 1'b1, 1'b0};
2159: data_out = {8'd109, 8'd221, 1'b1, 1'b0};
2160: data_out = {8'd145, 8'd221, 1'b1, 1'b0};
2161: data_out = {8'd168, 8'd221, 1'b1, 1'b0};
2162: data_out = {8'd169, 8'd221, 1'b1, 1'b0};
2163: data_out = {8'd86, 8'd222, 1'b1, 1'b0};
2164: data_out = {8'd87, 8'd222, 1'b1, 1'b0};
2165: data_out = {8'd108, 8'd222, 1'b1, 1'b0};
2166: data_out = {8'd109, 8'd222, 1'b1, 1'b0};
2167: data_out = {8'd145, 8'd222, 1'b1, 1'b0};
2168: data_out = {8'd146, 8'd222, 1'b1, 1'b0};
2169: data_out = {8'd167, 8'd222, 1'b1, 1'b0};
2170: data_out = {8'd168, 8'd222, 1'b1, 1'b0};
2171: data_out = {8'd87, 8'd223, 1'b1, 1'b0};
2172: data_out = {8'd108, 8'd223, 1'b1, 1'b0};
2173: data_out = {8'd146, 8'd223, 1'b1, 1'b0};
2174: data_out = {8'd167, 8'd223, 1'b1, 1'b0};
2175: data_out = {8'd87, 8'd224, 1'b1, 1'b0};
2176: data_out = {8'd88, 8'd224, 1'b1, 1'b0};
2177: data_out = {8'd107, 8'd224, 1'b1, 1'b0};
2178: data_out = {8'd108, 8'd224, 1'b1, 1'b0};
2179: data_out = {8'd146, 8'd224, 1'b1, 1'b0};
2180: data_out = {8'd147, 8'd224, 1'b1, 1'b0};
2181: data_out = {8'd166, 8'd224, 1'b1, 1'b0};
2182: data_out = {8'd167, 8'd224, 1'b1, 1'b0};
2183: data_out = {8'd88, 8'd225, 1'b1, 1'b0};
2184: data_out = {8'd89, 8'd225, 1'b1, 1'b0};
2185: data_out = {8'd107, 8'd225, 1'b1, 1'b0};
2186: data_out = {8'd147, 8'd225, 1'b1, 1'b0};
2187: data_out = {8'd165, 8'd225, 1'b1, 1'b0};
2188: data_out = {8'd166, 8'd225, 1'b1, 1'b0};
2189: data_out = {8'd89, 8'd226, 1'b1, 1'b0};
2190: data_out = {8'd90, 8'd226, 1'b1, 1'b0};
2191: data_out = {8'd106, 8'd226, 1'b1, 1'b0};
2192: data_out = {8'd107, 8'd226, 1'b1, 1'b0};
2193: data_out = {8'd147, 8'd226, 1'b1, 1'b0};
2194: data_out = {8'd148, 8'd226, 1'b1, 1'b0};
2195: data_out = {8'd164, 8'd226, 1'b1, 1'b0};
2196: data_out = {8'd165, 8'd226, 1'b1, 1'b0};
2197: data_out = {8'd90, 8'd227, 1'b1, 1'b0};
2198: data_out = {8'd91, 8'd227, 1'b1, 1'b0};
2199: data_out = {8'd105, 8'd227, 1'b1, 1'b0};
2200: data_out = {8'd106, 8'd227, 1'b1, 1'b0};
2201: data_out = {8'd148, 8'd227, 1'b1, 1'b0};
2202: data_out = {8'd149, 8'd227, 1'b1, 1'b0};
2203: data_out = {8'd163, 8'd227, 1'b1, 1'b0};
2204: data_out = {8'd164, 8'd227, 1'b1, 1'b0};
2205: data_out = {8'd91, 8'd228, 1'b1, 1'b0};
2206: data_out = {8'd92, 8'd228, 1'b1, 1'b0};
2207: data_out = {8'd105, 8'd228, 1'b1, 1'b0};
2208: data_out = {8'd149, 8'd228, 1'b1, 1'b0};
2209: data_out = {8'd162, 8'd228, 1'b1, 1'b0};
2210: data_out = {8'd163, 8'd228, 1'b1, 1'b0};
2211: data_out = {8'd92, 8'd229, 1'b1, 1'b0};
2212: data_out = {8'd93, 8'd229, 1'b1, 1'b0};
2213: data_out = {8'd104, 8'd229, 1'b1, 1'b0};
2214: data_out = {8'd105, 8'd229, 1'b1, 1'b0};
2215: data_out = {8'd149, 8'd229, 1'b1, 1'b0};
2216: data_out = {8'd150, 8'd229, 1'b1, 1'b0};
2217: data_out = {8'd161, 8'd229, 1'b1, 1'b0};
2218: data_out = {8'd162, 8'd229, 1'b1, 1'b0};
2219: data_out = {8'd93, 8'd230, 1'b1, 1'b0};
2220: data_out = {8'd94, 8'd230, 1'b1, 1'b0};
2221: data_out = {8'd104, 8'd230, 1'b1, 1'b0};
2222: data_out = {8'd150, 8'd230, 1'b1, 1'b0};
2223: data_out = {8'd160, 8'd230, 1'b1, 1'b0};
2224: data_out = {8'd161, 8'd230, 1'b1, 1'b0};
2225: data_out = {8'd94, 8'd231, 1'b1, 1'b0};
2226: data_out = {8'd95, 8'd231, 1'b1, 1'b0};
2227: data_out = {8'd96, 8'd231, 1'b1, 1'b0};
2228: data_out = {8'd103, 8'd231, 1'b1, 1'b0};
2229: data_out = {8'd104, 8'd231, 1'b1, 1'b0};
2230: data_out = {8'd150, 8'd231, 1'b1, 1'b0};
2231: data_out = {8'd151, 8'd231, 1'b1, 1'b0};
2232: data_out = {8'd158, 8'd231, 1'b1, 1'b0};
2233: data_out = {8'd159, 8'd231, 1'b1, 1'b0};
2234: data_out = {8'd160, 8'd231, 1'b1, 1'b0};
2235: data_out = {8'd96, 8'd232, 1'b1, 1'b0};
2236: data_out = {8'd97, 8'd232, 1'b1, 1'b0};
2237: data_out = {8'd103, 8'd232, 1'b1, 1'b0};
2238: data_out = {8'd151, 8'd232, 1'b1, 1'b0};
2239: data_out = {8'd157, 8'd232, 1'b1, 1'b0};
2240: data_out = {8'd158, 8'd232, 1'b1, 1'b0};
2241: data_out = {8'd97, 8'd233, 1'b1, 1'b0};
2242: data_out = {8'd98, 8'd233, 1'b1, 1'b0};
2243: data_out = {8'd102, 8'd233, 1'b1, 1'b0};
2244: data_out = {8'd103, 8'd233, 1'b1, 1'b0};
2245: data_out = {8'd151, 8'd233, 1'b1, 1'b0};
2246: data_out = {8'd152, 8'd233, 1'b1, 1'b0};
2247: data_out = {8'd156, 8'd233, 1'b1, 1'b0};
2248: data_out = {8'd157, 8'd233, 1'b1, 1'b0};
2249: data_out = {8'd98, 8'd234, 1'b1, 1'b0};
2250: data_out = {8'd99, 8'd234, 1'b1, 1'b0};
2251: data_out = {8'd100, 8'd234, 1'b1, 1'b0};
2252: data_out = {8'd101, 8'd234, 1'b1, 1'b0};
2253: data_out = {8'd102, 8'd234, 1'b1, 1'b0};
2254: data_out = {8'd152, 8'd234, 1'b1, 1'b0};
2255: data_out = {8'd153, 8'd234, 1'b1, 1'b0};
2256: data_out = {8'd154, 8'd234, 1'b1, 1'b0};
2257: data_out = {8'd155, 8'd234, 1'b1, 1'b0};
2258: data_out = {8'd156, 8'd234, 1'b1, 1'b0};
2259: data_out = {8'd100, 8'd235, 1'b1, 1'b0};
2260: data_out = {8'd101, 8'd235, 1'b1, 1'b0};
2261: data_out = {8'd153, 8'd235, 1'b1, 1'b0};
2262: data_out = {8'd154, 8'd235, 1'b1, 1'b1};




            default: data_out = '0;
        endcase
    end

endmodule
