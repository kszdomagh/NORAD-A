//////////////////////////////////////////////////////////////////////////////
/*
 Module name:   vector_pkg
 Author:        kszdom
 Description:  module used for holding all constants for vector stuff
 */
//////////////////////////////////////////////////////////////////////////////
package vector_pkg;

    // Parameters for 8 bit DAC vector output;
    localparam DAC_WIDTH = 8;
    localparam OUT_WIDTH = DAC_WIDTH;

    localparam Y_D0 = 7;
    localparam Y_D1 = 6;
    localparam Y_D2 = 5;
    localparam Y_D3 = 4;
    localparam Y_D4 = 3;
    localparam Y_D5 = 2;
    localparam Y_D6 = 1;
    localparam Y_D7 = 8;

    localparam X_D0 = 7;
    localparam X_D1 = 6;
    localparam X_D2 = 5;
    localparam X_D3 = 4;
    localparam X_D4 = 3;
    localparam X_D5 = 2;
    localparam X_D6 = 1;
    localparam X_D7 = 8;


    //PARAMETERS FOR VECTOR DISPLAY 255x255
    localparam VECTOR_MAX = 255;
    localparam VECTOR_MIN = 0;

    localparam CEASE_CYCLES = 2;



    //PARAMETERS FOR DATA
    localparam ADDRESSWIDTH = 16;
    localparam DATAWIDTH = 18;

endpackage
