//////////////////////////////////////////////////////////////////////////////
/*
 Module name:   ROM_pkg
 Author:        kszdom
 Description:  module used for holding all constants related to images in ROM memory
 */
//////////////////////////////////////////////////////////////////////////////
package ROM_pkg;

    // START OF ADRESSES FOR ROM IMAGES
    localparam ADR_MAP_START = 0;

    localparam ADR_FRAME_START = 42;

    localparam ADR_CURSOR_START = 48;



endpackage
